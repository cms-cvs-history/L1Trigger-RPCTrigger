-- Wed Oct 19 17:37:15 2005
library ieee;
use ieee.std_logic_1164.all;
use work.std_logic_1164_ktp.all;
use work.RPC_PAC_def.all;

package RPC_PAC_patt is

constant TT_EPACS_COUNT		:natural := 12; 
constant TT_TPACS_COUNT		:natural := 0; 
constant TT_REF_GROUP_NUMBERS	:natural := 1;
constant TT_GBSORT_INPUTS	:natural := 12; 

constant PACLogPlainsDecl	:TPACLogPlainsDecl := (
  --PAC_INDEX
  --|   PAC_MODEL
  --|   |      logplain 1 size .........logplain 6 size
   (0,  E, (  72,  56,   8,  40,  40,  24))
  ,(1,  E, (  72,  56,   8,  40,  40,  24))
  ,(2,  E, (  72,  56,   8,  40,  40,  24))
  ,(3,  E, (  72,  56,   8,  40,  40,  24))
  ,(4,  E, (  72,  56,   8,  40,  40,  24))
  ,(5,  E, (  72,  56,   8,  40,  40,  24))
  ,(6,  E, (  72,  56,   8,  40,  40,  24))
  ,(7,  E, (  72,  56,   8,  40,  40,  24))
  ,(8,  E, (  72,  56,   8,  40,  40,  24))
  ,(9,  E, (  72,  56,   8,  40,  40,  24))
  ,(10, E, (  72,  56,   8,  40,  40,  24))
  ,(11, E, (  72,  56,   8,  40,  40,  24))
  
);

constant LogPlainConn		:TLogPlainConn := (
  --PAC_INDEX   Logplane        LinkChannel     LinkLeftBit
  --| PAC_MODEL |       Link    |       LogPlaneLeftBit
  --|      |    |       |       |       |       |       LinkBitsCount
  --------------------------------------------------------------
   (0,    E,    0,      0,      0,      0,       0,      72) 
  ,(0,    E,    1,      1,      0,      0,       0,      56) 
  ,(0,    E,    2,      2,      0,      0,       0,       8) 
  ,(0,    E,    3,      3,      0,      0,       0,      40) 
  ,(0,    E,    4,      4,      0,      0,       0,      40) 
  ,(0,    E,    5,      5,      0,      0,       0,      24)  
  ,(0,    E,    0,      6,      0,      0,       0,      72) 
  ,(0,    E,    1,      7,      0,      0,       0,      56) 
  ,(0,    E,    2,      8,      0,      0,       0,       8) 
  ,(0,    E,    3,      9,      0,      0,       0,      40) 
  ,(0,    E,    4,     10,      0,      0,       0,      40) 
  ,(0,    E,    5,     11,      0,      0,       0,      24)  
  
  ,(1,    E,    0,      0,      0,      0,       8,      72) 
  ,(1,    E,    1,      1,      0,      0,       8,      56) 
  ,(1,    E,    2,      2,      0,      0,       8,       8) 
  ,(1,    E,    3,      3,      0,      0,       8,      40) 
  ,(1,    E,    4,      4,      0,      0,       8,      40) 
  ,(1,    E,    5,      5,      0,      0,       8,      24) 	 
  ,(1,    E,    0,      6,      0,      0,       8,      72)  
  ,(1,    E,    1,      7,      0,      0,       8,      56)  
  ,(1,    E,    2,      8,      0,      0,       8,       8)  
  ,(1,    E,    3,      9,      0,      0,       8,      40)  
  ,(1,    E,    4,     10,      0,      0,       8,      40)  
  ,(1,    E,    5,     11,      0,      0,       8,      24) 	
 
  ,(2,    E,    0,      0,      0,      0,      16,      72) 
  ,(2,    E,    1,      1,      0,      0,      16,      56) 
  ,(2,    E,    2,      2,      0,      0,      16,       8) 
  ,(2,    E,    3,      3,      0,      0,      16,      40) 
  ,(2,    E,    4,      4,      0,      0,      16,      40) 
  ,(2,    E,    5,      5,      0,      0,      16,      24) 
  ,(2,    E,    0,      6,      0,      0,      16,      72) 
  ,(2,    E,    1,      7,      0,      0,      16,      56) 
  ,(2,    E,    2,      8,      0,      0,      16,       8) 
  ,(2,    E,    3,      9,      0,      0,      16,      40) 
  ,(2,    E,    4,     10,      0,      0,      16,      40) 
  ,(2,    E,    5,     11,      0,      0,      16,      24) 
  
  ,(3,    E,    0,      0,      0,      0,      24,      72)
  ,(3,    E,    1,      1,      0,      0,      24,      56) 
  ,(3,    E,    2,      2,      0,      0,      24,       8) 
  ,(3,    E,    3,      3,      0,      0,      24,      40) 
  ,(3,    E,    4,      4,      0,      0,      24,      40) 
  ,(3,    E,    5,      5,      0,      0,      24,      24)  
  ,(3,    E,    0,      6,      0,      0,      24,      72)
  ,(3,    E,    1,      7,      0,      0,      24,      56) 
  ,(3,    E,    2,      8,      0,      0,      24,       8) 
  ,(3,    E,    3,      9,      0,      0,      24,      40) 
  ,(3,    E,    4,     10,      0,      0,      24,      40) 
  ,(3,    E,    5,     11,      0,      0,      24,      24)  
  
  ,(4,    E,    0,      0,      0,      0,      32,      64)  
  ,(4,    E,    0,      0,      1,     64,       0,       8)
  ,(4,    E,    1,      1,      0,      0,      32,      56)
  ,(4,    E,    2,      2,      0,      0,      32,       8)
  ,(4,    E,    3,      3,      0,      0,      32,      40)
  ,(4,    E,    4,      4,      0,      0,      32,      40)
  ,(4,    E,    5,      5,      0,      0,      32,      24)
  ,(4,    E,    0,      6,      0,      0,      32,      64)  
  ,(4,    E,    0,      6,      1,     64,       0,       8)
  ,(4,    E,    1,      7,      0,      0,      32,      56)
  ,(4,    E,    2,      8,      0,      0,      32,       8)
  ,(4,    E,    3,      9,      0,      0,      32,      40)
  ,(4,    E,    4,     10,      0,      0,      32,      40)
  ,(4,    E,    5,     11,      0,      0,      32,      24)

  ,(5,    E,    0,      0,      0,      0,      40,      56)
  ,(5,    E,    0,      0,      1,     56,       0,      16)
  ,(5,    E,    1,      1,      0,      0,      40,      56)
  ,(5,    E,    2,      2,      0,      0,      40,       8)
  ,(5,    E,    3,      3,      0,      0,      40,      40)
  ,(5,    E,    4,      4,      0,      0,      40,      40)
  ,(5,    E,    5,      5,      0,      0,      40,      24)
  ,(5,    E,    0,      6,      0,      0,      40,      56)
  ,(5,    E,    0,      6,      1,     56,       0,      16)
  ,(5,    E,    1,      7,      0,      0,      40,      56)
  ,(5,    E,    2,      8,      0,      0,      40,       8)
  ,(5,    E,    3,      9,      0,      0,      40,      40)
  ,(5,    E,    4,     10,      0,      0,      40,      40)
  ,(5,    E,    5,     11,      0,      0,      40,      24)
  
  ,(6,    E,    0,      0,      0,      0,      48,      48)
  ,(6,    E,    0,      0,      1,     48,       0,      24)
  ,(6,    E,    1,      1,      0,      0,      48,      48)     
  ,(6,    E,    1,      1,      1,     48,       0,       8)
  ,(6,    E,    2,      2,      0,      0,      48,       8)
  ,(6,    E,    3,      3,      0,      0,      48,      40)
  ,(6,    E,    4,      4,      0,      0,      48,      40)
  ,(6,    E,    5,      5,      0,      0,      48,      24)
  ,(6,    E,    0,      6,      0,      0,      48,      48)
  ,(6,    E,    0,      6,      1,     48,       0,      24)
  ,(6,    E,    1,      7,      0,      0,      48,      48)     
  ,(6,    E,    1,      7,      1,     48,       0,       8)
  ,(6,    E,    2,      8,      0,      0,      48,       8)
  ,(6,    E,    3,      9,      0,      0,      48,      40)
  ,(6,    E,    4,     10,      0,      0,      48,      40)
  ,(6,    E,    5,     11,      0,      0,      48,      24)
  
  ,(7,    E,    0,      0,      0,      0,      56,      40)
  ,(7,    E,    0,      0,      1,     40,       0,      32)
  ,(7,    E,    1,      1,      0,      0,      56,      40)
  ,(7,    E,    1,      1,      1,     40,       0,      16)
  ,(7,    E,    2,      2,      0,      0,      56,       8)
  ,(7,    E,    3,      3,      0,      0,      56,      40)
  ,(7,    E,    4,      4,      0,      0,      56,      40)
  ,(7,    E,    5,      5,      0,      0,      56,      24)
  ,(7,    E,    0,      6,      0,      0,      56,      40)
  ,(7,    E,    0,      6,      1,     40,       0,      32)
  ,(7,    E,    1,      7,      0,      0,      56,      40)
  ,(7,    E,    1,      7,      1,     40,       0,      16)
  ,(7,    E,    2,      8,      0,      0,      56,       8)
  ,(7,    E,    3,      9,      0,      0,      56,      40)
  ,(7,    E,    4,     10,      0,      0,      56,      40)
  ,(7,    E,    5,     11,      0,      0,      56,      24)

  ,(8,    E,    0,      0,      0,      0,      64,      32)
  ,(8,    E,    0,      0,      1,     32,       0,      40)
  ,(8,    E,    1,      1,      0,      0,      64,      32)
  ,(8,    E,    1,      1,      1,     32,       0,      24)
  ,(8,    E,    2,      2,      0,      0,      64,       8)
  ,(8,    E,    3,      3,      0,      0,      64,      32)
  ,(8,    E,    3,      3,      1,     32,       0,       8)  
  ,(8,    E,    4,      4,      0,      0,      64,      32)
  ,(8,    E,    4,      4,      1,     32,       0,       8)  
  ,(8,    E,    5,      5,      0,      0,      64,      24)
  ,(8,    E,    0,      6,      0,      0,      64,      32)
  ,(8,    E,    0,      6,      1,     32,       0,      40)
  ,(8,    E,    1,      7,      0,      0,      64,      32)
  ,(8,    E,    1,      7,      1,     32,       0,      24)
  ,(8,    E,    2,      8,      0,      0,      64,       8)
  ,(8,    E,    3,      9,      0,      0,      64,      32)
  ,(8,    E,    3,      9,      1,     32,       0,       8)  
  ,(8,    E,    4,     10,      0,      0,      64,      32)
  ,(8,    E,    4,     10,      1,     32,       0,       8)  
  ,(8,    E,    5,     11,      0,      0,      64,      24)

  ,(9,    E,    0,      0,      0,      0,      72,      24)
  ,(9,    E,    0,      0,      1,     24,       0,      48)
  ,(9,    E,    1,      1,      0,      0,      72,      24)
  ,(9,    E,    1,      1,      1,     24,       0,      32)
  ,(9,    E,    2,      2,      0,      0,      72,       8)
  ,(9,    E,    3,      3,      0,      0,      72,      24)
  ,(9,    E,    3,      3,      1,     24,       0,      16)
  ,(9,    E,    4,      4,      0,      0,      72,      24)
  ,(9,    E,    4,      4,      1,     24,       0,      16)
  ,(9,    E,    5,      5,      0,      0,      72,      24)
  ,(9,    E,    0,      6,      0,      0,      72,      24)
  ,(9,    E,    0,      6,      1,     24,       0,      48)
  ,(9,    E,    1,      7,      0,      0,      72,      24)
  ,(9,    E,    1,      7,      1,     24,       0,      32)
  ,(9,    E,    2,      8,      0,      0,      72,       8)
  ,(9,    E,    3,      9,      0,      0,      72,      24)
  ,(9,    E,    3,      9,      1,     24,       0,      16)
  ,(9,    E,    4,     10,      0,      0,      72,      24)
  ,(9,    E,    4,     10,      1,     24,       0,      16)
  ,(9,    E,    5,     11,      0,      0,      72,      24)

  ,(10,   E,    0,      0,      0,      0,      80,      16)
  ,(10,   E,    0,      0,      1,     16,       0,      56)
  ,(10,   E,    1,      1,      0,      0,      80,      16)
  ,(10,   E,    1,      1,      1,     16,       0,      40)
  ,(10,   E,    2,      2,      0,      0,      80,       8)
  ,(10,   E,    3,      3,      0,      0,      80,      16)
  ,(10,   E,    3,      3,      1,     16,       0,      24)
  ,(10,   E,    4,      4,      0,      0,      80,      16)
  ,(10,   E,    4,      4,      1,     16,       0,      24)
  ,(10,   E,    5,      5,      0,      0,      80,      16)
  ,(10,   E,    5,      5,      1,     16,       0,       8)
  ,(10,   E,    0,      6,      0,      0,      80,      16)
  ,(10,   E,    0,      6,      1,     16,       0,      56)
  ,(10,   E,    1,      7,      0,      0,      80,      16)
  ,(10,   E,    1,      7,      1,     16,       0,      40)
  ,(10,   E,    2,      8,      0,      0,      80,       8)
  ,(10,   E,    3,      9,      0,      0,      80,      16)
  ,(10,   E,    3,      9,      1,     16,       0,      24)
  ,(10,   E,    4,     10,      0,      0,      80,      16)
  ,(10,   E,    4,     10,      1,     16,       0,      24)
  ,(10,   E,    5,     11,      0,      0,      80,      16)
  ,(10,   E,    5,     11,      1,     16,       0,       8)

  ,(11,   E,    0,      0,      0,      0,      88,       8)
  ,(11,   E,    0,      0,      1,      8,       0,      64)
  ,(11,   E,    1,      1,      0,      0,      88,       8)
  ,(11,   E,    1,      1,      1,      8,       0,      48)
  ,(11,   E,    2,      2,      0,      0,      88,       8)
  ,(11,   E,    3,      3,      0,      0,      88,       8)
  ,(11,   E,    3,      3,      1,      8,       0,      32)
  ,(11,   E,    4,      4,      0,      0,      88,       8)
  ,(11,   E,    4,      4,      1,      8,       0,      32)
  ,(11,   E,    5,      5,      0,      0,      88,       8)
  ,(11,   E,    5,      5,      0,      8,       0,      16)  
  ,(11,   E,    0,      6,      0,      0,      88,       8)
  ,(11,   E,    0,      6,      1,      8,       0,      64)
  ,(11,   E,    1,      7,      0,      0,      88,       8)
  ,(11,   E,    1,      7,      1,      8,       0,      48)
  ,(11,   E,    2,      8,      0,      0,      88,       8)
  ,(11,   E,    3,      9,      0,      0,      88,       8)
  ,(11,   E,    3,      9,      1,      8,       0,      32)
  ,(11,   E,    4,     10,      0,      0,      88,       8)
  ,(11,   E,    4,     10,      1,      8,       0,      32)
  ,(11,   E,    5,     11,      0,      0,      88,       8)
  ,(11,   E,    5,     11,      0,      8,       0,      16)  

);

constant GBSortDecl		:TGBSortDecl := (  
  --PAC_INDEX
  --|   PAC_MODEL
  --|	 |   GBSORT_INPUT_INDEX			
   (0,   E,  0)
	,(1,   E,  1)
	,(2,   E,  2)
	,(3,   E,  3)
	,(4,   E,  4)
	,(5,   E,  5)	
	,(6,   E,  6)
	,(7,   E,  7)
	,(8,   E,  8)
	,(9,   E,  9)
	,(10,  E,  10)      
	,(11,  E,  11)
);
constant PACCellQuality :TPACCellQuality := (
--   654321
 (0,"001111",1), 
 (0,"010111",1), 
 (0,"011011",1), 
 (0,"011101",1), 
 (0,"011110",1), 
 (0,"011111",2), 
 (0,"100111",1), 
 (0,"101011",1), 
 (0,"101101",1), 
 (0,"101110",1), 
 (0,"101111",2), 
 (0,"110011",1), 
 (0,"110101",1), 
 (0,"110110",1), 
 (0,"110111",2), 
 (0,"111001",1), 
 (0,"111010",1), 
 (0,"111011",2), 
 (0,"111100",1), 
 (0,"111101",2), 
 (0,"111110",2), 
 (0,"111111",3), 
 (1,"000111",0), 
 (1,"001011",0), 
 (1,"001101",0), 
 (1,"001110",0), 
 (1,"001111",1)
);
constant PACPattTable :TPACPattTable := (
--PAC_INDEX
--| PAC_MODEL
--| | Ref Group Index
--| | | Qualit Tab index
--| | | |  Plane1  Plane2  Plane3  Plane4  Plane5  Plane6  sign code  pat number
 ( 0, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 31) -- 0
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 31) -- 1
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 31) -- 2
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 31) -- 3
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 31) -- 4
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 31) -- 5
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 31) -- 6
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 31) -- 7
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 8
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 9
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 10
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 11
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 12
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 13
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 14
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 15
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 31) -- 16
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 31) -- 17
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 31) -- 18
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 31) -- 19
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 31) -- 20
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 31) -- 21
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 31) -- 22
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 31) -- 23
,( 0, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 24
,( 0, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 25
,( 0, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 26
,( 0, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 27
,( 0, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 28
,( 0, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 29
,( 0, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 30
,( 0, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 31
,( 0, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 31) -- 32
,( 0, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),(10,10)), 1, 31) -- 33
,( 0, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(11,11)), 1, 31) -- 34
,( 0, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(12,12)), 1, 31) -- 35
,( 0, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(13,13)), 1, 31) -- 36
,( 0, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(14,14)), 1, 31) -- 37
,( 0, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(15,15)), 1, 31) -- 38
,( 0, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(16,16)), 1, 31) -- 39
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 31) -- 40
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 1, 31) -- 41
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 1, 31) -- 42
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 1, 31) -- 43
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 1, 31) -- 44
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 1, 31) -- 45
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 1, 31) -- 46
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 1, 31) -- 47
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 31) -- 48
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 31) -- 49
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(17,17),(10,10)), 1, 31) -- 50
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(18,18),(11,11)), 1, 31) -- 51
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(19,19),(12,12)), 1, 31) -- 52
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(20,20),(13,13)), 1, 31) -- 53
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(21,21),(14,14)), 1, 31) -- 54
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(22,22),(15,15)), 1, 31) -- 55
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 31) -- 56
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 31) -- 57
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 31) -- 58
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 31) -- 59
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 31) -- 60
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 31) -- 61
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 31) -- 62
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 31) -- 63
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 30) -- 64
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 30) -- 65
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 30) -- 66
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 30) -- 67
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 30) -- 68
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 30) -- 69
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 30) -- 70
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 30) -- 71
,( 0, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 29) -- 72
,( 0, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 29) -- 73
,( 0, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(17,17),(10,10)), 1, 29) -- 74
,( 0, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(18,18),(11,11)), 1, 29) -- 75
,( 0, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(19,19),(12,12)), 1, 29) -- 76
,( 0, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(20,20),(13,13)), 1, 29) -- 77
,( 0, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(21,21),(14,14)), 1, 29) -- 78
,( 0, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(22,22),(15,15)), 1, 29) -- 79
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 27) -- 80
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 27) -- 81
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),(10,10)), 1, 27) -- 82
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(11,11)), 1, 27) -- 83
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(12,12)), 1, 27) -- 84
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(13,13)), 1, 27) -- 85
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(14,14)), 1, 27) -- 86
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(15,15)), 1, 27) -- 87
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 25) -- 88
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 25) -- 89
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 25) -- 90
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 25) -- 91
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 25) -- 92
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 25) -- 93
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 25) -- 94
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 25) -- 95
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 25) -- 96
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 25) -- 97
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),(10,10)), 1, 25) -- 98
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(11,11)), 1, 25) -- 99
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(12,12)), 1, 25) -- 100
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(13,13)), 1, 25) -- 101
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(14,14)), 1, 25) -- 102
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(15,15)), 1, 25) -- 103
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 104
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 105
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 106
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 107
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 108
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 109
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 110
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 111
,( 0, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 112
,( 0, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 113
,( 0, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 114
,( 0, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 115
,( 0, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 116
,( 0, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 117
,( 0, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 118
,( 0, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 119
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 22) -- 120
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 22) -- 121
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 22) -- 122
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(17,17),(10,10)), 1, 22) -- 123
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(18,18),(11,11)), 1, 22) -- 124
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(19,19),(12,12)), 1, 22) -- 125
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(20,20),(13,13)), 1, 22) -- 126
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(21,21),(14,14)), 1, 22) -- 127
,( 0, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 22) -- 128
,( 0, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 22) -- 129
,( 0, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 22) -- 130
,( 0, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),(10,10)), 1, 22) -- 131
,( 0, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(11,11)), 1, 22) -- 132
,( 0, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(12,12)), 1, 22) -- 133
,( 0, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(13,13)), 1, 22) -- 134
,( 0, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(14,14)), 1, 22) -- 135
,( 0, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 21) -- 136
,( 0, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 21) -- 137
,( 0, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 21) -- 138
,( 0, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 21) -- 139
,( 0, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 21) -- 140
,( 0, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 21) -- 141
,( 0, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 21) -- 142
,( 0, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 21) -- 143
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 21) -- 144
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 21) -- 145
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 21) -- 146
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 21) -- 147
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 21) -- 148
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 21) -- 149
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 21) -- 150
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 21) -- 151
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 21) -- 152
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 21) -- 153
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 21) -- 154
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 21) -- 155
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 21) -- 156
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 21) -- 157
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 21) -- 158
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 21) -- 159
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 20) -- 160
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 20) -- 161
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 20) -- 162
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 20) -- 163
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 20) -- 164
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 20) -- 165
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 20) -- 166
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 20) -- 167
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 168
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 169
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 170
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 171
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 172
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 173
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 174
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 175
,( 0, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 20) -- 176
,( 0, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 20) -- 177
,( 0, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 20) -- 178
,( 0, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 20) -- 179
,( 0, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 20) -- 180
,( 0, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 20) -- 181
,( 0, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 20) -- 182
,( 0, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 20) -- 183
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 19) -- 184
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 19) -- 185
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 19) -- 186
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 19) -- 187
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 19) -- 188
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 19) -- 189
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 19) -- 190
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 19) -- 191
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 19) -- 192
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 19) -- 193
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 19) -- 194
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 19) -- 195
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 19) -- 196
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 19) -- 197
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 19) -- 198
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 19) -- 199
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 19) -- 200
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 19) -- 201
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),(10,10)), 1, 19) -- 202
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(11,11)), 1, 19) -- 203
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(12,12)), 1, 19) -- 204
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(13,13)), 1, 19) -- 205
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(14,14)), 1, 19) -- 206
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(15,15)), 1, 19) -- 207
,( 0, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 208
,( 0, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 209
,( 0, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 210
,( 0, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 211
,( 0, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 212
,( 0, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 213
,( 0, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 214
,( 0, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 215
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 216
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 217
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 218
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 219
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 220
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 221
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 222
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 223
,( 0, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 224
,( 0, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 225
,( 0, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 226
,( 0, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 227
,( 0, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 228
,( 0, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 229
,( 0, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 230
,( 0, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 231
,( 0, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 232
,( 0, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 233
,( 0, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 234
,( 0, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 235
,( 0, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 236
,( 0, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 237
,( 0, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 238
,( 0, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 239
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 18) -- 240
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 18) -- 241
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 18) -- 242
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 18) -- 243
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 18) -- 244
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 18) -- 245
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 18) -- 246
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 18) -- 247
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 248
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 249
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 250
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 251
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 252
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 253
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 254
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 255
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 256
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 257
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 258
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 259
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 260
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 261
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 262
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 263
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 17) -- 264
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 17) -- 265
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 17) -- 266
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 17) -- 267
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 17) -- 268
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 17) -- 269
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 17) -- 270
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 17) -- 271
,( 0, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 17) -- 272
,( 0, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 17) -- 273
,( 0, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 17) -- 274
,( 0, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),(10,10)), 1, 17) -- 275
,( 0, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),(11,11)), 1, 17) -- 276
,( 0, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(12,12)), 1, 17) -- 277
,( 0, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(13,13)), 1, 17) -- 278
,( 0, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(14,14)), 1, 17) -- 279
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 280
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 281
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 282
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 283
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 284
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 285
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 286
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 287
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 17) -- 288
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 17) -- 289
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 17) -- 290
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),(10,10)), 1, 17) -- 291
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(11,11)), 1, 17) -- 292
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(12,12)), 1, 17) -- 293
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(13,13)), 1, 17) -- 294
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(14,14)), 1, 17) -- 295
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(13,13),( 6, 6)), 1, 17) -- 296
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(14,14),( 7, 7)), 1, 17) -- 297
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(15,15),( 8, 8)), 1, 17) -- 298
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(16,16),( 9, 9)), 1, 17) -- 299
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(17,17),(10,10)), 1, 17) -- 300
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(18,18),(11,11)), 1, 17) -- 301
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(19,19),(12,12)), 1, 17) -- 302
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(20,20),(13,13)), 1, 17) -- 303
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 17) -- 304
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 17) -- 305
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 17) -- 306
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 17) -- 307
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 17) -- 308
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(18,18),(10,10)), 1, 17) -- 309
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(19,19),(11,11)), 1, 17) -- 310
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(20,20),(12,12)), 1, 17) -- 311
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 16) -- 312
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 16) -- 313
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 16) -- 314
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 16) -- 315
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 16) -- 316
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(18,18),(10,10)), 1, 16) -- 317
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(19,19),(11,11)), 1, 16) -- 318
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(20,20),(12,12)), 1, 16) -- 319
,( 0, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 16) -- 320
,( 0, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 16) -- 321
,( 0, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 16) -- 322
,( 0, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 16) -- 323
,( 0, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 16) -- 324
,( 0, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 16) -- 325
,( 0, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 16) -- 326
,( 0, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 16) -- 327
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 328
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 329
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 330
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 331
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 332
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 333
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 334
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 335
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 336
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 337
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 338
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 339
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 340
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 341
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 342
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 343
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(13,13),( 6, 6)), 1, 15) -- 344
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(14,14),( 7, 7)), 1, 15) -- 345
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(15,15),( 8, 8)), 1, 15) -- 346
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(16,16),( 9, 9)), 1, 15) -- 347
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(17,17),(10,10)), 1, 15) -- 348
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(18,18),(11,11)), 1, 15) -- 349
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(19,19),(12,12)), 1, 15) -- 350
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(20,20),(13,13)), 1, 15) -- 351
,( 0, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 352
,( 0, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 353
,( 0, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 354
,( 0, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 355
,( 0, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 356
,( 0, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 357
,( 0, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 358
,( 0, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 359
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 6, 6)), 1, 15) -- 360
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 7, 7)), 1, 15) -- 361
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 8, 8)), 1, 15) -- 362
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 9, 9)), 1, 15) -- 363
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),(10,10)), 1, 15) -- 364
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(11,11)), 1, 15) -- 365
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(12,12)), 1, 15) -- 366
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(13,13)), 1, 15) -- 367
,( 0, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 368
,( 0, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 369
,( 0, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 370
,( 0, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 371
,( 0, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 372
,( 0, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 373
,( 0, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 374
,( 0, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 375
,( 0, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 15) -- 376
,( 0, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 15) -- 377
,( 0, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 15) -- 378
,( 0, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 15) -- 379
,( 0, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 15) -- 380
,( 0, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(18,18),(10,10)), 1, 15) -- 381
,( 0, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(19,19),(11,11)), 1, 15) -- 382
,( 0, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(20,20),(12,12)), 1, 15) -- 383
,( 0, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 384
,( 0, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 385
,( 0, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 386
,( 0, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 387
,( 0, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 388
,( 0, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 389
,( 0, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 390
,( 0, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 391
,( 0, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 392
,( 0, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 393
,( 0, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 394
,( 0, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 395
,( 0, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 396
,( 0, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 397
,( 0, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 398
,( 0, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 399
,( 0, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 400
,( 0, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 401
,( 0, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 402
,( 0, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 403
,( 0, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 404
,( 0, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 405
,( 0, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 406
,( 0, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 407
,( 0, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 6, 6)), 1, 15) -- 408
,( 0, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 7, 7)), 1, 15) -- 409
,( 0, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 8, 8)), 1, 15) -- 410
,( 0, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 9, 9)), 1, 15) -- 411
,( 0, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),(10,10)), 1, 15) -- 412
,( 0, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(11,11)), 1, 15) -- 413
,( 0, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(12,12)), 1, 15) -- 414
,( 0, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(13,13)), 1, 15) -- 415
,( 0, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 416
,( 0, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 417
,( 0, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 418
,( 0, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 419
,( 0, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 420
,( 0, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 421
,( 0, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 422
,( 0, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 423
,( 0, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 424
,( 0, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 425
,( 0, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 426
,( 0, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 427
,( 0, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 428
,( 0, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 429
,( 0, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 430
,( 0, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 431
,( 0, E,0,0,((36,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 432
,( 0, E,0,0,((38,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 433
,( 0, E,0,0,((40,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 434
,( 0, E,0,0,((42,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 435
,( 0, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 4, 7)), 1, 13) -- 436
,( 0, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 6, 9)), 1, 13) -- 437
,( 0, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),( 8,11)), 1, 13) -- 438
,( 0, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),(10,13)), 1, 13) -- 439
,( 0, E,0,0,((36,39),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 13) -- 440
,( 0, E,0,0,((38,41),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 13) -- 441
,( 0, E,0,0,((40,43),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 13) -- 442
,( 0, E,0,0,((42,45),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 13) -- 443
,( 0, E,0,0,((36,39),(28,28),( 1, 1),(15,15),(14,14),( 4, 7)), 1, 13) -- 444
,( 0, E,0,0,((38,41),(30,30),( 3, 3),(17,17),(16,16),( 6, 9)), 1, 13) -- 445
,( 0, E,0,0,((40,43),(32,32),( 5, 5),(19,19),(18,18),( 8,11)), 1, 13) -- 446
,( 0, E,0,0,((42,45),(34,34),( 7, 7),(21,21),(20,20),(10,13)), 1, 13) -- 447
,( 0, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 4, 7)), 1, 12) -- 448
,( 0, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 6, 9)), 1, 12) -- 449
,( 0, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 8,11)), 1, 12) -- 450
,( 0, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(10,13)), 1, 12) -- 451
,( 0, E,0,0,((36,39),(26,27),( 0, 1),(14,14),(11,11),( 0, 3)), 1, 12) -- 452
,( 0, E,0,0,((38,41),(28,29),( 2, 3),(16,16),(13,13),( 2, 5)), 1, 12) -- 453
,( 0, E,0,0,((40,43),(30,31),( 4, 5),(18,18),(15,15),( 4, 7)), 1, 12) -- 454
,( 0, E,0,0,((42,45),(32,33),( 6, 7),(20,20),(17,17),( 6, 9)), 1, 12) -- 455
,( 0, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(10,11),( 2, 5)), 1, 12) -- 456
,( 0, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(12,13),( 4, 7)), 1, 12) -- 457
,( 0, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(14,15),( 6, 9)), 1, 12) -- 458
,( 0, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(16,17),( 8,11)), 1, 12) -- 459
,( 0, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 12) -- 460
,( 0, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),( 8,11)), 1, 12) -- 461
,( 0, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),(10,13)), 1, 12) -- 462
,( 0, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(12,15)), 1, 12) -- 463
,( 0, E,0,0,((38,41),(28,29),( 0, 1),(14,14),(10,11),( 2, 5)), 1, 11) -- 464
,( 0, E,0,0,((40,43),(30,31),( 2, 3),(16,16),(12,13),( 4, 7)), 1, 11) -- 465
,( 0, E,0,0,((42,45),(32,33),( 4, 5),(18,18),(14,15),( 6, 9)), 1, 11) -- 466
,( 0, E,0,0,((44,47),(34,35),( 6, 7),(20,20),(16,17),( 8,11)), 1, 11) -- 467
,( 0, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 11) -- 468
,( 0, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 11) -- 469
,( 0, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 11) -- 470
,( 0, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 11) -- 471
,( 0, E,0,0,((40,41),(28,29),( 0, 1),(14,15),(12,12),( 2, 3)), 1, 11) -- 472
,( 0, E,0,0,((42,43),(30,31),( 2, 3),(16,17),(14,14),( 4, 5)), 1, 11) -- 473
,( 0, E,0,0,((44,45),(32,33),( 4, 5),(18,19),(16,16),( 6, 7)), 1, 11) -- 474
,( 0, E,0,0,((46,47),(34,35),( 6, 7),(20,21),(18,18),( 8, 9)), 1, 11) -- 475
,( 0, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 476
,( 0, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 477
,( 0, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(10,13)), 1, 11) -- 478
,( 0, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(12,15)), 1, 11) -- 479
,( 0, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,12),( 4, 7)), 1, 11) -- 480
,( 0, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,14),( 6, 9)), 1, 11) -- 481
,( 0, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,16),( 8,11)), 1, 11) -- 482
,( 0, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,18),(10,13)), 1, 11) -- 483
,( 0, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(10,11),( 4, 7)), 1, 10) -- 484
,( 0, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(12,13),( 6, 9)), 1, 10) -- 485
,( 0, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(14,15),( 8,11)), 1, 10) -- 486
,( 0, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(16,17),(10,13)), 1, 10) -- 487
,( 0, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(12,13),( 4, 7)), 1, 10) -- 488
,( 0, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(14,15),( 6, 9)), 1, 10) -- 489
,( 0, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(16,17),( 8,11)), 1, 10) -- 490
,( 0, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(18,19),(10,13)), 1, 10) -- 491
,( 0, E,0,0,((40,43),(30,31),( 1, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 492
,( 0, E,0,0,((42,45),(32,33),( 3, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 493
,( 0, E,0,0,((44,47),(34,35),( 5, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 494
,( 0, E,0,0,((46,49),(36,37),( 7, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 495
,( 0, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 8,11)), 1, 10) -- 496
,( 0, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),(10,13)), 1, 10) -- 497
,( 0, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(12,15)), 1, 10) -- 498
,( 0, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(14,17)), 1, 10) -- 499
,( 0, E,0,0,((40,43),(28,29),( 0, 0),(12,13),( 8, 9),( 0, 3)), 1, 10) -- 500
,( 0, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(10,11),( 2, 5)), 1, 10) -- 501
,( 0, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(12,13),( 4, 7)), 1, 10) -- 502
,( 0, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(14,15),( 6, 9)), 1, 10) -- 503
,( 0, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,12),( 4, 7)), 1, 10) -- 504
,( 0, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,14),( 6, 9)), 1, 10) -- 505
,( 0, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,16),( 8,11)), 1, 10) -- 506
,( 0, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,18),(10,13)), 1, 10) -- 507
,( 0, E,0,0,((42,43),(30,30),( 0, 1),(13,13),(10,11),( 0, 3)), 1, 10) -- 508
,( 0, E,0,0,((44,45),(32,32),( 2, 3),(15,15),(12,13),( 2, 5)), 1, 10) -- 509
,( 0, E,0,0,((46,47),(34,34),( 4, 5),(17,17),(14,15),( 4, 7)), 1, 10) -- 510
,( 0, E,0,0,((48,49),(36,36),( 6, 7),(19,19),(16,17),( 6, 9)), 1, 10) -- 511
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 512
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 513
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 514
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 515
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),( 6, 9)), 1,  9) -- 516
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),( 8,11)), 1,  9) -- 517
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(10,13)), 1,  9) -- 518
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(12,15)), 1,  9) -- 519
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 2, 5)), 1,  9) -- 520
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 4, 7)), 1,  9) -- 521
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 6, 9)), 1,  9) -- 522
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 8,11)), 1,  9) -- 523
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(10,11),( 4, 7)), 1,  9) -- 524
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(12,13),( 6, 9)), 1,  9) -- 525
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(14,15),( 8,11)), 1,  9) -- 526
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(16,17),(10,13)), 1,  9) -- 527
,( 0, E,0,0,((40,43),(29,29),( 0, 0),(12,13),(10,11),( 4, 7)), 1,  9) -- 528
,( 0, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(12,13),( 6, 9)), 1,  9) -- 529
,( 0, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(14,15),( 8,11)), 1,  9) -- 530
,( 0, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(16,17),(10,13)), 1,  9) -- 531
,( 0, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),( 8,11)), 1,  9) -- 532
,( 0, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),(10,13)), 1,  9) -- 533
,( 0, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(12,15)), 1,  9) -- 534
,( 0, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(14,17)), 1,  9) -- 535
,( 0, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(14,15),( 8,11)), 1,  9) -- 536
,( 0, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(16,17),(10,13)), 1,  9) -- 537
,( 0, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(18,19),(12,15)), 1,  9) -- 538
,( 0, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(20,21),(14,17)), 1,  9) -- 539
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),(10,13)), 1,  9) -- 540
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(12,15)), 1,  9) -- 541
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(14,17)), 1,  9) -- 542
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(16,19)), 1,  9) -- 543
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 1)), 1,  9) -- 544
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 3)), 1,  9) -- 545
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 5)), 1,  9) -- 546
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 7)), 1,  9) -- 547
,( 0, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 8,11)), 1,  9) -- 548
,( 0, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),(10,13)), 1,  9) -- 549
,( 0, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(12,15)), 1,  9) -- 550
,( 0, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(14,17)), 1,  9) -- 551
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(13,13),(10,11),( 8,11)), 1,  9) -- 552
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(15,15),(12,13),(10,13)), 1,  9) -- 553
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(17,17),(14,15),(12,15)), 1,  9) -- 554
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(19,19),(16,17),(14,17)), 1,  9) -- 555
,( 0, E,0,0,((42,42),(29,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1,  9) -- 556
,( 0, E,0,0,((44,44),(31,31),( 2, 3),(16,17),(14,15),( 8,11)), 1,  9) -- 557
,( 0, E,0,0,((46,46),(33,33),( 4, 5),(18,19),(16,17),(10,13)), 1,  9) -- 558
,( 0, E,0,0,((48,48),(35,35),( 6, 7),(20,21),(18,19),(12,15)), 1,  9) -- 559
,( 0, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(11,11),( 6, 9)), 1,  9) -- 560
,( 0, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(13,13),( 8,11)), 1,  9) -- 561
,( 0, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(15,15),(10,13)), 1,  9) -- 562
,( 0, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(17,17),(12,15)), 1,  9) -- 563
,( 0, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 0, 3)), 1,  9) -- 564
,( 0, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 2, 5)), 1,  9) -- 565
,( 0, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 4, 7)), 1,  9) -- 566
,( 0, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),( 6, 9)), 1,  9) -- 567
,( 0, E,0,0,((40,41),(29,29),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 568
,( 0, E,0,0,((42,43),(31,31),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 569
,( 0, E,0,0,((44,45),(33,33),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 570
,( 0, E,0,0,((46,47),(35,35),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 571
,( 0, E,0,0,((46,49),(32,33),( 0, 1),(12,13),( 8, 9),( 6, 6)), 1,  9) -- 572
,( 0, E,0,0,((48,51),(34,35),( 2, 3),(14,15),(10,11),( 8, 8)), 1,  9) -- 573
,( 0, E,0,0,((50,53),(36,37),( 4, 5),(16,17),(12,13),(10,10)), 1,  9) -- 574
,( 0, E,0,0,((52,55),(38,39),( 6, 7),(18,19),(14,15),(12,12)), 1,  9) -- 575
,( 0, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),(10,13)), 1,  9) -- 576
,( 0, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(12,15)), 1,  9) -- 577
,( 0, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(14,17)), 1,  9) -- 578
,( 0, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(16,19)), 1,  9) -- 579
,( 0, E,0,0,((40,43),(29,29),( 0, 1),(13,13),(10,11),( 0, 3)), 1,  9) -- 580
,( 0, E,0,0,((42,45),(31,31),( 2, 3),(15,15),(12,13),( 2, 5)), 1,  9) -- 581
,( 0, E,0,0,((44,47),(33,33),( 4, 5),(17,17),(14,15),( 4, 7)), 1,  9) -- 582
,( 0, E,0,0,((46,49),(35,35),( 6, 7),(19,19),(16,17),( 6, 9)), 1,  9) -- 583
,( 0, E,0,0,((44,47),(32,33),( 1, 1),(13,13),(10,11),( 4, 4)), 1,  9) -- 584
,( 0, E,0,0,((46,49),(34,35),( 3, 3),(15,15),(12,13),( 6, 6)), 1,  9) -- 585
,( 0, E,0,0,((48,51),(36,37),( 5, 5),(17,17),(14,15),( 8, 8)), 1,  9) -- 586
,( 0, E,0,0,((50,53),(38,39),( 7, 7),(19,19),(16,17),(10,10)), 1,  9) -- 587
,( 0, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(10,13),( 6, 9)), 1,  8) -- 588
,( 0, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(12,15),( 8,11)), 1,  8) -- 589
,( 0, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(14,17),(10,13)), 1,  8) -- 590
,( 0, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(16,19),(12,15)), 1,  8) -- 591
,( 0, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 6, 9),( 6, 9)), 1,  8) -- 592
,( 0, E,0,0,((46,49),(32,35),( 2, 3),(12,15),( 8,11),( 8,11)), 1,  8) -- 593
,( 0, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(10,13),(10,13)), 1,  8) -- 594
,( 0, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(12,15),(12,15)), 1,  8) -- 595
,( 0, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 596
,( 0, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 597
,( 0, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 598
,( 0, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 599
,( 0, E,0,0,((48,51),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 600
,( 0, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 601
,( 0, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 602
,( 0, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 603
,( 0, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  7) -- 604
,( 0, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  7) -- 605
,( 0, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  7) -- 606
,( 0, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  7) -- 607
,( 0, E,0,1,((48,51),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 608
,( 0, E,0,1,((50,53),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 609
,( 0, E,0,1,((52,55),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 610
,( 0, E,0,1,((54,57),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 611
,( 0, E,0,1,((48,51),(32,35),( 0, 1),(14,17),(99,99),(99,99)), 1,  7) -- 612
,( 0, E,0,1,((50,53),(34,37),( 2, 3),(16,19),(99,99),(99,99)), 1,  7) -- 613
,( 0, E,0,1,((52,55),(36,39),( 4, 5),(18,21),(99,99),(99,99)), 1,  7) -- 614
,( 0, E,0,1,((54,57),(38,41),( 6, 7),(20,23),(99,99),(99,99)), 1,  7) -- 615
,( 0, E,0,1,((44,47),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 616
,( 0, E,0,1,((46,49),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 617
,( 0, E,0,1,((48,51),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 618
,( 0, E,0,1,((50,53),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 619
,( 0, E,0,1,((52,55),(34,37),( 0, 1),(10,13),(99,99),(99,99)), 1,  6) -- 620
,( 0, E,0,1,((54,57),(36,39),( 2, 3),(12,15),(99,99),(99,99)), 1,  6) -- 621
,( 0, E,0,1,((56,59),(38,41),( 4, 5),(14,17),(99,99),(99,99)), 1,  6) -- 622
,( 0, E,0,1,((58,61),(40,43),( 6, 7),(16,19),(99,99),(99,99)), 1,  6) -- 623
,( 0, E,0,1,((46,49),(31,31),( 0, 0),(14,15),(99,99),(99,99)), 1,  5) -- 624
,( 0, E,0,1,((48,51),(33,33),( 2, 2),(16,17),(99,99),(99,99)), 1,  5) -- 625
,( 0, E,0,1,((50,53),(35,35),( 4, 4),(18,19),(99,99),(99,99)), 1,  5) -- 626
,( 0, E,0,1,((52,55),(37,37),( 6, 6),(20,21),(99,99),(99,99)), 1,  5) -- 627
,( 0, E,0,1,((42,45),(28,31),( 0, 1),(20,23),(99,99),(99,99)), 1,  5) -- 628
,( 0, E,0,1,((44,47),(30,33),( 2, 3),(22,25),(99,99),(99,99)), 1,  5) -- 629
,( 0, E,0,1,((46,49),(32,35),( 4, 5),(24,27),(99,99),(99,99)), 1,  5) -- 630
,( 0, E,0,1,((48,51),(34,37),( 6, 7),(26,29),(99,99),(99,99)), 1,  5) -- 631
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 632
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 633
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 634
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 635
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 636
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 637
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 638
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 639
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 0, 31) -- 640
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 0, 31) -- 641
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 0, 31) -- 642
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 0, 31) -- 643
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 0, 31) -- 644
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 0, 31) -- 645
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 0, 31) -- 646
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 0, 31) -- 647
,( 0, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 648
,( 0, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 649
,( 0, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 650
,( 0, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 651
,( 0, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 652
,( 0, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 653
,( 0, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 654
,( 0, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 655
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 656
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 657
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 658
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 659
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 660
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 661
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 662
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 663
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 664
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 665
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 666
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 667
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 668
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 669
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 670
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 671
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 672
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 673
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 674
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 675
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 676
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 677
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 678
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 679
,( 0, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(15,15),( 8, 8)), 0, 31) -- 680
,( 0, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(16,16),( 9, 9)), 0, 31) -- 681
,( 0, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(17,17),(10,10)), 0, 31) -- 682
,( 0, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(18,18),(11,11)), 0, 31) -- 683
,( 0, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(19,19),(12,12)), 0, 31) -- 684
,( 0, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(20,20),(13,13)), 0, 31) -- 685
,( 0, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(21,21),(14,14)), 0, 31) -- 686
,( 0, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(22,22),(15,15)), 0, 31) -- 687
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 29) -- 688
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),(10,10)), 0, 29) -- 689
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(11,11)), 0, 29) -- 690
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(12,12)), 0, 29) -- 691
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(13,13)), 0, 29) -- 692
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(14,14)), 0, 29) -- 693
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(15,15)), 0, 29) -- 694
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(16,16)), 0, 29) -- 695
,( 0, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 28) -- 696
,( 0, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 28) -- 697
,( 0, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 28) -- 698
,( 0, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 28) -- 699
,( 0, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 28) -- 700
,( 0, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 28) -- 701
,( 0, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 28) -- 702
,( 0, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 28) -- 703
,( 0, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 26) -- 704
,( 0, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 26) -- 705
,( 0, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 26) -- 706
,( 0, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 26) -- 707
,( 0, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 26) -- 708
,( 0, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 26) -- 709
,( 0, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 26) -- 710
,( 0, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 26) -- 711
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 25) -- 712
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 25) -- 713
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 25) -- 714
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 25) -- 715
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 25) -- 716
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 25) -- 717
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 25) -- 718
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 25) -- 719
,( 0, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 25) -- 720
,( 0, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 25) -- 721
,( 0, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 25) -- 722
,( 0, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 25) -- 723
,( 0, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 25) -- 724
,( 0, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 25) -- 725
,( 0, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 25) -- 726
,( 0, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 25) -- 727
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 25) -- 728
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 25) -- 729
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 25) -- 730
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 25) -- 731
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 25) -- 732
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 25) -- 733
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 25) -- 734
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 25) -- 735
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 24) -- 736
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 24) -- 737
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 24) -- 738
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 24) -- 739
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 24) -- 740
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 24) -- 741
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 24) -- 742
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 24) -- 743
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 23) -- 744
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 23) -- 745
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 23) -- 746
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 23) -- 747
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 23) -- 748
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 23) -- 749
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 23) -- 750
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 23) -- 751
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 22) -- 752
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 22) -- 753
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 22) -- 754
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 22) -- 755
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 22) -- 756
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 22) -- 757
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 22) -- 758
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 22) -- 759
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 22) -- 760
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 22) -- 761
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 22) -- 762
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 22) -- 763
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 22) -- 764
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 22) -- 765
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 22) -- 766
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 22) -- 767
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 768
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 769
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 770
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 771
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 772
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 773
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 774
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 775
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 20) -- 776
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 20) -- 777
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 20) -- 778
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 20) -- 779
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 20) -- 780
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 20) -- 781
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 20) -- 782
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 20) -- 783
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),(10,10)), 0, 20) -- 784
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(11,11)), 0, 20) -- 785
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(12,12)), 0, 20) -- 786
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(13,13)), 0, 20) -- 787
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(14,14)), 0, 20) -- 788
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(15,15)), 0, 20) -- 789
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(16,16)), 0, 20) -- 790
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(17,17)), 0, 20) -- 791
,( 0, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 792
,( 0, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 793
,( 0, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 794
,( 0, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 795
,( 0, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 796
,( 0, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 797
,( 0, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 798
,( 0, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 799
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(11,11)), 0, 19) -- 800
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(12,12)), 0, 19) -- 801
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(13,13)), 0, 19) -- 802
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(14,14)), 0, 19) -- 803
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(15,15)), 0, 19) -- 804
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(16,16)), 0, 19) -- 805
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(17,17)), 0, 19) -- 806
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(18,18)), 0, 19) -- 807
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 808
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 809
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 810
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 811
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 812
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 813
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 814
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 815
,( 0, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(17,17),(10,10)), 0, 19) -- 816
,( 0, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(18,18),(11,11)), 0, 19) -- 817
,( 0, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(19,19),(12,12)), 0, 19) -- 818
,( 0, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(20,20),(13,13)), 0, 19) -- 819
,( 0, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(21,21),(14,14)), 0, 19) -- 820
,( 0, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(22,22),(15,15)), 0, 19) -- 821
,( 0, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(23,23),(16,16)), 0, 19) -- 822
,( 0, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(24,24),(17,17)), 0, 19) -- 823
,( 0, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 824
,( 0, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 825
,( 0, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 826
,( 0, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 827
,( 0, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 828
,( 0, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 829
,( 0, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 830
,( 0, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 831
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(17,17),(10,10)), 0, 18) -- 832
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(18,18),(11,11)), 0, 18) -- 833
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(19,19),(12,12)), 0, 18) -- 834
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(20,20),(13,13)), 0, 18) -- 835
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(21,21),(14,14)), 0, 18) -- 836
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(22,22),(15,15)), 0, 18) -- 837
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(23,23),(16,16)), 0, 18) -- 838
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(24,24),(17,17)), 0, 18) -- 839
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 840
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 841
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 842
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 843
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 844
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 845
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 846
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 847
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 18) -- 848
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 18) -- 849
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 18) -- 850
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 18) -- 851
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 18) -- 852
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 18) -- 853
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 18) -- 854
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 18) -- 855
,( 0, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(17,17),(10,10)), 0, 18) -- 856
,( 0, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(18,18),(11,11)), 0, 18) -- 857
,( 0, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(19,19),(12,12)), 0, 18) -- 858
,( 0, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(20,20),(13,13)), 0, 18) -- 859
,( 0, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(21,21),(14,14)), 0, 18) -- 860
,( 0, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(22,22),(15,15)), 0, 18) -- 861
,( 0, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(23,23),(16,16)), 0, 18) -- 862
,( 0, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(24,24),(17,17)), 0, 18) -- 863
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 18) -- 864
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 18) -- 865
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 18) -- 866
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 18) -- 867
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 18) -- 868
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 18) -- 869
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 18) -- 870
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 18) -- 871
,( 0, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 872
,( 0, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 873
,( 0, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 874
,( 0, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 875
,( 0, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 876
,( 0, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 877
,( 0, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 878
,( 0, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 879
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(11,11)), 0, 18) -- 880
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(12,12)), 0, 18) -- 881
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(13,13)), 0, 18) -- 882
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(14,14)), 0, 18) -- 883
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(15,15)), 0, 18) -- 884
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(16,16)), 0, 18) -- 885
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(17,17)), 0, 18) -- 886
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(18,18)), 0, 18) -- 887
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 888
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 889
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 890
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 891
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 892
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 893
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 894
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 895
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(17,17),(11,11)), 0, 17) -- 896
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(18,18),(12,12)), 0, 17) -- 897
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(19,19),(13,13)), 0, 17) -- 898
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(20,20),(14,14)), 0, 17) -- 899
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(21,21),(15,15)), 0, 17) -- 900
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(22,22),(16,16)), 0, 17) -- 901
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(23,23),(17,17)), 0, 17) -- 902
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(24,24),(18,18)), 0, 17) -- 903
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 904
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 905
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 906
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 907
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 908
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 909
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 910
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 911
,( 0, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 912
,( 0, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 913
,( 0, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 914
,( 0, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 915
,( 0, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 916
,( 0, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 917
,( 0, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 918
,( 0, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 919
,( 0, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(11,11)), 0, 17) -- 920
,( 0, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(12,12)), 0, 17) -- 921
,( 0, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(13,13)), 0, 17) -- 922
,( 0, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(14,14)), 0, 17) -- 923
,( 0, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(15,15)), 0, 17) -- 924
,( 0, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(16,16)), 0, 17) -- 925
,( 0, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(17,17)), 0, 17) -- 926
,( 0, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(18,18)), 0, 17) -- 927
,( 0, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 17) -- 928
,( 0, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 17) -- 929
,( 0, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 17) -- 930
,( 0, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 17) -- 931
,( 0, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 17) -- 932
,( 0, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 17) -- 933
,( 0, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 17) -- 934
,( 0, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 17) -- 935
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 16) -- 936
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 16) -- 937
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 16) -- 938
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 16) -- 939
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 16) -- 940
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 16) -- 941
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 16) -- 942
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 16) -- 943
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(12,12)), 0, 16) -- 944
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(13,13)), 0, 16) -- 945
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(14,14)), 0, 16) -- 946
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(15,15)), 0, 16) -- 947
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(16,16)), 0, 16) -- 948
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(17,17)), 0, 16) -- 949
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(18,18)), 0, 16) -- 950
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(19,19)), 0, 16) -- 951
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 952
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 953
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 954
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 955
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 956
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 957
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 958
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 959
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 16) -- 960
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 16) -- 961
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 16) -- 962
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 16) -- 963
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 16) -- 964
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 16) -- 965
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 16) -- 966
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 16) -- 967
,( 0, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(17,17),(10,10)), 0, 16) -- 968
,( 0, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(18,18),(11,11)), 0, 16) -- 969
,( 0, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(19,19),(12,12)), 0, 16) -- 970
,( 0, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(20,20),(13,13)), 0, 16) -- 971
,( 0, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(21,21),(14,14)), 0, 16) -- 972
,( 0, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(22,22),(15,15)), 0, 16) -- 973
,( 0, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(23,23),(16,16)), 0, 16) -- 974
,( 0, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(24,24),(17,17)), 0, 16) -- 975
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(11,11)), 0, 16) -- 976
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(12,12)), 0, 16) -- 977
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(13,13)), 0, 16) -- 978
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(14,14)), 0, 16) -- 979
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(15,15)), 0, 16) -- 980
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(16,16)), 0, 16) -- 981
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(17,17)), 0, 16) -- 982
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(18,18)), 0, 16) -- 983
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 984
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 985
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 986
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 987
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 988
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 989
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 990
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 991
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(12,12)), 0, 15) -- 992
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(13,13)), 0, 15) -- 993
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(14,14)), 0, 15) -- 994
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(15,15)), 0, 15) -- 995
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(16,16)), 0, 15) -- 996
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(17,17)), 0, 15) -- 997
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(18,18)), 0, 15) -- 998
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(19,19)), 0, 15) -- 999
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(12,12)), 0, 15) -- 1000
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(13,13)), 0, 15) -- 1001
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(14,14)), 0, 15) -- 1002
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(15,15)), 0, 15) -- 1003
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(16,16)), 0, 15) -- 1004
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(17,17)), 0, 15) -- 1005
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(18,18)), 0, 15) -- 1006
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(19,19)), 0, 15) -- 1007
,( 0, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 15) -- 1008
,( 0, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 15) -- 1009
,( 0, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 15) -- 1010
,( 0, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 15) -- 1011
,( 0, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 15) -- 1012
,( 0, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 15) -- 1013
,( 0, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 15) -- 1014
,( 0, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 15) -- 1015
,( 0, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 1016
,( 0, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 1017
,( 0, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 1018
,( 0, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 1019
,( 0, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 1020
,( 0, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 1021
,( 0, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 1022
,( 0, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 1023
,( 0, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 1024
,( 0, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 1025
,( 0, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 1026
,( 0, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 1027
,( 0, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(20,21),(12,15)), 0, 14) -- 1028
,( 0, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(22,23),(14,17)), 0, 14) -- 1029
,( 0, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(24,25),(16,19)), 0, 14) -- 1030
,( 0, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(26,27),(18,21)), 0, 14) -- 1031
,( 0, E,0,0,((28,31),(22,23),( 0, 1),(18,18),(18,19),(10,13)), 0, 14) -- 1032
,( 0, E,0,0,((30,33),(24,25),( 2, 3),(20,20),(20,21),(12,15)), 0, 14) -- 1033
,( 0, E,0,0,((32,35),(26,27),( 4, 5),(22,22),(22,23),(14,17)), 0, 14) -- 1034
,( 0, E,0,0,((34,37),(28,29),( 6, 7),(24,24),(24,25),(16,19)), 0, 14) -- 1035
,( 0, E,0,0,((26,27),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 13) -- 1036
,( 0, E,0,0,((28,29),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 13) -- 1037
,( 0, E,0,0,((30,31),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 13) -- 1038
,( 0, E,0,0,((32,33),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 13) -- 1039
,( 0, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 1040
,( 0, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 1041
,( 0, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 1042
,( 0, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 1043
,( 0, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(18,19),(10,13)), 0, 12) -- 1044
,( 0, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(20,21),(12,15)), 0, 12) -- 1045
,( 0, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(22,23),(14,17)), 0, 12) -- 1046
,( 0, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(24,25),(16,19)), 0, 12) -- 1047
,( 0, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,20),(12,15)), 0, 12) -- 1048
,( 0, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,22),(14,17)), 0, 12) -- 1049
,( 0, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,24),(16,19)), 0, 12) -- 1050
,( 0, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,26),(18,21)), 0, 12) -- 1051
,( 0, E,0,0,((24,25),(20,21),( 0, 0),(17,17),(18,19),(10,13)), 0, 12) -- 1052
,( 0, E,0,0,((26,27),(22,23),( 2, 2),(19,19),(20,21),(12,15)), 0, 12) -- 1053
,( 0, E,0,0,((28,29),(24,25),( 4, 4),(21,21),(22,23),(14,17)), 0, 12) -- 1054
,( 0, E,0,0,((30,31),(26,27),( 6, 6),(23,23),(24,25),(16,19)), 0, 12) -- 1055
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 1056
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 1057
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 1058
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 1059
,( 0, E,0,0,((24,27),(20,21),( 0, 1),(18,18),(19,19),(10,13)), 0, 11) -- 1060
,( 0, E,0,0,((26,29),(22,23),( 2, 3),(20,20),(21,21),(12,15)), 0, 11) -- 1061
,( 0, E,0,0,((28,31),(24,25),( 4, 5),(22,22),(23,23),(14,17)), 0, 11) -- 1062
,( 0, E,0,0,((30,33),(26,27),( 6, 7),(24,24),(25,25),(16,19)), 0, 11) -- 1063
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),(10,13)), 0, 11) -- 1064
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),(12,15)), 0, 11) -- 1065
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(14,17)), 0, 11) -- 1066
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(16,19)), 0, 11) -- 1067
,( 0, E,0,0,((24,27),(20,21),( 0, 0),(16,17),(18,19),( 6, 9)), 0, 11) -- 1068
,( 0, E,0,0,((26,29),(22,23),( 2, 2),(18,19),(20,21),( 8,11)), 0, 11) -- 1069
,( 0, E,0,0,((28,31),(24,25),( 4, 4),(20,21),(22,23),(10,13)), 0, 11) -- 1070
,( 0, E,0,0,((30,33),(26,27),( 6, 6),(22,23),(24,25),(12,15)), 0, 11) -- 1071
,( 0, E,0,0,((24,27),(22,23),( 1, 1),(18,19),(20,21),(10,13)), 0, 11) -- 1072
,( 0, E,0,0,((26,29),(24,25),( 3, 3),(20,21),(22,23),(12,15)), 0, 11) -- 1073
,( 0, E,0,0,((28,31),(26,27),( 5, 5),(22,23),(24,25),(14,17)), 0, 11) -- 1074
,( 0, E,0,0,((30,33),(28,29),( 7, 7),(24,25),(26,27),(16,19)), 0, 11) -- 1075
,( 0, E,0,0,((24,27),(22,22),( 1, 1),(19,19),(22,23),(14,17)), 0, 11) -- 1076
,( 0, E,0,0,((26,29),(24,24),( 3, 3),(21,21),(24,25),(16,19)), 0, 11) -- 1077
,( 0, E,0,0,((28,31),(26,26),( 5, 5),(23,23),(26,27),(18,21)), 0, 11) -- 1078
,( 0, E,0,0,((30,33),(28,28),( 7, 7),(25,25),(28,29),(20,23)), 0, 11) -- 1079
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,18),(21,21),(14,17)), 0, 11) -- 1080
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,20),(23,23),(16,19)), 0, 11) -- 1081
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,22),(25,25),(18,21)), 0, 11) -- 1082
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,24),(27,27),(20,23)), 0, 11) -- 1083
,( 0, E,0,0,((20,23),(19,19),( 0, 1),(18,19),(20,21),(12,15)), 0, 10) -- 1084
,( 0, E,0,0,((22,25),(21,21),( 2, 3),(20,21),(22,23),(14,17)), 0, 10) -- 1085
,( 0, E,0,0,((24,27),(23,23),( 4, 5),(22,23),(24,25),(16,19)), 0, 10) -- 1086
,( 0, E,0,0,((26,29),(25,25),( 6, 7),(24,25),(26,27),(18,21)), 0, 10) -- 1087
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(19,19),(22,22),(10,13)), 0, 10) -- 1088
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(21,21),(24,24),(12,15)), 0, 10) -- 1089
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(23,23),(26,26),(14,17)), 0, 10) -- 1090
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(25,25),(28,28),(16,19)), 0, 10) -- 1091
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 6, 9)), 0, 10) -- 1092
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 8,11)), 0, 10) -- 1093
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),(10,13)), 0, 10) -- 1094
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),(12,15)), 0, 10) -- 1095
,( 0, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(14,17)), 0, 10) -- 1096
,( 0, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(16,19)), 0, 10) -- 1097
,( 0, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(18,21)), 0, 10) -- 1098
,( 0, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(20,23)), 0, 10) -- 1099
,( 0, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(22,23),(14,17)), 0, 10) -- 1100
,( 0, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(24,25),(16,19)), 0, 10) -- 1101
,( 0, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(26,27),(18,21)), 0, 10) -- 1102
,( 0, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(28,29),(20,23)), 0, 10) -- 1103
,( 0, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(20,21),( 8,11)), 0, 10) -- 1104
,( 0, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(22,23),(10,13)), 0, 10) -- 1105
,( 0, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(24,25),(12,15)), 0, 10) -- 1106
,( 0, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(26,27),(14,17)), 0, 10) -- 1107
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,20),( 6, 9)), 0, 10) -- 1108
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,22),( 8,11)), 0, 10) -- 1109
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,24),(10,13)), 0, 10) -- 1110
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,26),(12,15)), 0, 10) -- 1111
,( 0, E,0,0,((23,23),(20,20),( 0, 0),(17,17),(18,19),( 6, 9)), 0, 10) -- 1112
,( 0, E,0,0,((25,25),(22,22),( 2, 2),(19,19),(20,21),( 8,11)), 0, 10) -- 1113
,( 0, E,0,0,((27,27),(24,24),( 4, 4),(21,21),(22,23),(10,13)), 0, 10) -- 1114
,( 0, E,0,0,((29,29),(26,26),( 6, 6),(23,23),(24,25),(12,15)), 0, 10) -- 1115
,( 0, E,0,0,((22,23),(19,19),( 0, 0),(17,17),(20,20),(10,13)), 0, 10) -- 1116
,( 0, E,0,0,((24,25),(21,21),( 2, 2),(19,19),(22,22),(12,15)), 0, 10) -- 1117
,( 0, E,0,0,((26,27),(23,23),( 4, 4),(21,21),(24,24),(14,17)), 0, 10) -- 1118
,( 0, E,0,0,((28,29),(25,25),( 6, 6),(23,23),(26,26),(16,19)), 0, 10) -- 1119
,( 0, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(20,20),(10,13)), 0, 10) -- 1120
,( 0, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(22,22),(12,15)), 0, 10) -- 1121
,( 0, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(24,24),(14,17)), 0, 10) -- 1122
,( 0, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(26,26),(16,19)), 0, 10) -- 1123
,( 0, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(10,13)), 0,  9) -- 1124
,( 0, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(12,15)), 0,  9) -- 1125
,( 0, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(14,17)), 0,  9) -- 1126
,( 0, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(16,19)), 0,  9) -- 1127
,( 0, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(18,19),( 6, 9)), 0,  9) -- 1128
,( 0, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(20,21),( 8,11)), 0,  9) -- 1129
,( 0, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(22,23),(10,13)), 0,  9) -- 1130
,( 0, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(24,25),(12,15)), 0,  9) -- 1131
,( 0, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 1132
,( 0, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 1133
,( 0, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 1134
,( 0, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 1135
,( 0, E,0,0,((20,23),(20,20),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 1136
,( 0, E,0,0,((22,25),(22,22),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 1137
,( 0, E,0,0,((24,27),(24,24),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 1138
,( 0, E,0,0,((26,29),(26,26),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 1139
,( 0, E,0,0,((18,21),(18,19),( 1, 1),(20,21),(22,23),( 8,11)), 0,  9) -- 1140
,( 0, E,0,0,((20,23),(20,21),( 3, 3),(22,23),(24,25),(10,13)), 0,  9) -- 1141
,( 0, E,0,0,((22,25),(22,23),( 5, 5),(24,25),(26,27),(12,15)), 0,  9) -- 1142
,( 0, E,0,0,((24,27),(24,25),( 7, 7),(26,27),(28,29),(14,17)), 0,  9) -- 1143
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(21,21),( 6, 9)), 0,  9) -- 1144
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(23,23),( 8,11)), 0,  9) -- 1145
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(25,25),(10,13)), 0,  9) -- 1146
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(27,27),(12,15)), 0,  9) -- 1147
,( 0, E,0,0,((18,21),(18,19),( 0, 1),(20,21),(24,25),(14,17)), 0,  9) -- 1148
,( 0, E,0,0,((20,23),(20,21),( 2, 3),(22,23),(26,27),(16,19)), 0,  9) -- 1149
,( 0, E,0,0,((22,25),(22,23),( 4, 5),(24,25),(28,29),(18,21)), 0,  9) -- 1150
,( 0, E,0,0,((24,27),(24,25),( 6, 7),(26,27),(30,31),(20,23)), 0,  9) -- 1151
,( 0, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(21,21),(10,13)), 0,  9) -- 1152
,( 0, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(23,23),(12,15)), 0,  9) -- 1153
,( 0, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(25,25),(14,17)), 0,  9) -- 1154
,( 0, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(27,27),(16,19)), 0,  9) -- 1155
,( 0, E,0,0,((20,23),(19,19),( 0, 0),(17,17),(18,19),( 6, 9)), 0,  9) -- 1156
,( 0, E,0,0,((22,25),(21,21),( 2, 2),(19,19),(20,21),( 8,11)), 0,  9) -- 1157
,( 0, E,0,0,((24,27),(23,23),( 4, 4),(21,21),(22,23),(10,13)), 0,  9) -- 1158
,( 0, E,0,0,((26,29),(25,25),( 6, 6),(23,23),(24,25),(12,15)), 0,  9) -- 1159
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 1160
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 1161
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 1162
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 1163
,( 0, E,0,0,((20,23),(19,19),( 1, 1),(19,19),(22,23),(14,17)), 0,  9) -- 1164
,( 0, E,0,0,((22,25),(21,21),( 3, 3),(21,21),(24,25),(16,19)), 0,  9) -- 1165
,( 0, E,0,0,((24,27),(23,23),( 5, 5),(23,23),(26,27),(18,21)), 0,  9) -- 1166
,( 0, E,0,0,((26,29),(25,25),( 7, 7),(25,25),(28,29),(20,23)), 0,  9) -- 1167
,( 0, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 1168
,( 0, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 1169
,( 0, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 1170
,( 0, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 1171
,( 0, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(22,23),(12,15)), 0,  9) -- 1172
,( 0, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(24,25),(14,17)), 0,  9) -- 1173
,( 0, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(26,27),(16,19)), 0,  9) -- 1174
,( 0, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(28,29),(18,21)), 0,  9) -- 1175
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(19,19),(20,21),( 2, 5)), 0,  9) -- 1176
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(21,21),(22,23),( 4, 7)), 0,  9) -- 1177
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(23,23),(24,25),( 6, 9)), 0,  9) -- 1178
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(25,25),(26,27),( 8,11)), 0,  9) -- 1179
,( 0, E,0,0,((16,19),(16,17),( 0, 0),(19,19),(22,23),(10,13)), 0,  9) -- 1180
,( 0, E,0,0,((18,21),(18,19),( 2, 2),(21,21),(24,25),(12,15)), 0,  9) -- 1181
,( 0, E,0,0,((20,23),(20,21),( 4, 4),(23,23),(26,27),(14,17)), 0,  9) -- 1182
,( 0, E,0,0,((22,25),(22,23),( 6, 6),(25,25),(28,29),(16,19)), 0,  9) -- 1183
,( 0, E,0,0,((18,21),(18,19),( 0, 1),(20,20),(20,21),( 6, 7)), 0,  9) -- 1184
,( 0, E,0,0,((20,23),(20,21),( 2, 3),(22,22),(22,23),( 8, 9)), 0,  9) -- 1185
,( 0, E,0,0,((22,25),(22,23),( 4, 5),(24,24),(24,25),(10,11)), 0,  9) -- 1186
,( 0, E,0,0,((24,27),(24,25),( 6, 7),(26,26),(26,27),(12,13)), 0,  9) -- 1187
,( 0, E,0,0,((18,21),(18,19),( 0, 1),(19,19),(22,23),( 8,11)), 0,  9) -- 1188
,( 0, E,0,0,((20,23),(20,21),( 2, 3),(21,21),(24,25),(10,13)), 0,  9) -- 1189
,( 0, E,0,0,((22,25),(22,23),( 4, 5),(23,23),(26,27),(12,15)), 0,  9) -- 1190
,( 0, E,0,0,((24,27),(24,25),( 6, 7),(25,25),(28,29),(14,17)), 0,  9) -- 1191
,( 0, E,0,0,((18,19),(17,17),( 0, 0),(18,19),(20,21),(10,10)), 0,  9) -- 1192
,( 0, E,0,0,((20,21),(19,19),( 2, 2),(20,21),(22,23),(12,12)), 0,  9) -- 1193
,( 0, E,0,0,((22,23),(21,21),( 4, 4),(22,23),(24,25),(14,14)), 0,  9) -- 1194
,( 0, E,0,0,((24,25),(23,23),( 6, 6),(24,25),(26,27),(16,16)), 0,  9) -- 1195
,( 0, E,0,0,((22,23),(20,21),( 1, 1),(20,20),(22,22),( 6, 9)), 0,  9) -- 1196
,( 0, E,0,0,((24,25),(22,23),( 3, 3),(22,22),(24,24),( 8,11)), 0,  9) -- 1197
,( 0, E,0,0,((26,27),(24,25),( 5, 5),(24,24),(26,26),(10,13)), 0,  9) -- 1198
,( 0, E,0,0,((28,29),(26,27),( 7, 7),(26,26),(28,28),(12,15)), 0,  9) -- 1199
,( 0, E,0,0,((22,25),(20,21),( 0, 1),(16,17),(16,17),( 2, 5)), 0,  9) -- 1200
,( 0, E,0,0,((24,27),(22,23),( 2, 3),(18,19),(18,19),( 4, 7)), 0,  9) -- 1201
,( 0, E,0,0,((26,29),(24,25),( 4, 5),(20,21),(20,21),( 6, 9)), 0,  9) -- 1202
,( 0, E,0,0,((28,31),(26,27),( 6, 7),(22,23),(22,23),( 8,11)), 0,  9) -- 1203
,( 0, E,0,0,((22,22),(19,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 1204
,( 0, E,0,0,((24,24),(21,21),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 1205
,( 0, E,0,0,((26,26),(23,23),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 1206
,( 0, E,0,0,((28,28),(25,25),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 1207
,( 0, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(22,25),(12,12)), 0,  8) -- 1208
,( 0, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(24,27),(14,14)), 0,  8) -- 1209
,( 0, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(26,29),(16,16)), 0,  8) -- 1210
,( 0, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(28,31),(18,18)), 0,  8) -- 1211
,( 0, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(18,21),( 8,11)), 0,  8) -- 1212
,( 0, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(20,23),(10,13)), 0,  8) -- 1213
,( 0, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(22,25),(12,15)), 0,  8) -- 1214
,( 0, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(24,27),(14,17)), 0,  8) -- 1215
,( 0, E,0,0,((20,23),(18,21),( 0, 1),(18,21),(18,21),( 4, 4)), 0,  8) -- 1216
,( 0, E,0,0,((22,25),(20,23),( 2, 3),(20,23),(20,23),( 6, 6)), 0,  8) -- 1217
,( 0, E,0,0,((24,27),(22,25),( 4, 5),(22,25),(22,25),( 8, 8)), 0,  8) -- 1218
,( 0, E,0,0,((26,29),(24,27),( 6, 7),(24,27),(24,27),(10,10)), 0,  8) -- 1219
,( 0, E,0,0,((18,21),(16,19),( 0, 1),(16,19),(16,19),(99,99)), 0,  8) -- 1220
,( 0, E,0,0,((20,23),(18,21),( 2, 3),(18,21),(18,21),(99,99)), 0,  8) -- 1221
,( 0, E,0,0,((22,25),(20,23),( 4, 5),(20,23),(20,23),(99,99)), 0,  8) -- 1222
,( 0, E,0,0,((24,27),(22,25),( 6, 7),(22,25),(22,25),(99,99)), 0,  8) -- 1223
,( 0, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 1224
,( 0, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 1225
,( 0, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 1226
,( 0, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 1227
,( 0, E,0,0,((12,15),(14,17),( 0, 1),(18,21),(20,23),(99,99)), 0,  7) -- 1228
,( 0, E,0,0,((14,17),(16,19),( 2, 3),(20,23),(22,25),(99,99)), 0,  7) -- 1229
,( 0, E,0,0,((16,19),(18,21),( 4, 5),(22,25),(24,27),(99,99)), 0,  7) -- 1230
,( 0, E,0,0,((18,21),(20,23),( 6, 7),(24,27),(26,29),(99,99)), 0,  7) -- 1231
,( 0, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 1232
,( 0, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 1233
,( 0, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 1234
,( 0, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 1235
,( 0, E,0,1,((14,17),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  7) -- 1236
,( 0, E,0,1,((16,19),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  7) -- 1237
,( 0, E,0,1,((18,21),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  7) -- 1238
,( 0, E,0,1,((20,23),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  7) -- 1239
,( 0, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 1240
,( 0, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 1241
,( 0, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 1242
,( 0, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 1243
,( 0, E,0,1,((10,13),(14,17),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 1244
,( 0, E,0,1,((12,15),(16,19),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 1245
,( 0, E,0,1,((14,17),(18,21),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 1246
,( 0, E,0,1,((16,19),(20,23),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 1247
,( 0, E,0,1,(( 8,11),(12,15),( 0, 1),(20,23),(99,99),(99,99)), 0,  6) -- 1248
,( 0, E,0,1,((10,13),(14,17),( 2, 3),(22,25),(99,99),(99,99)), 0,  6) -- 1249
,( 0, E,0,1,((12,15),(16,19),( 4, 5),(24,27),(99,99),(99,99)), 0,  6) -- 1250
,( 0, E,0,1,((14,17),(18,21),( 6, 7),(26,29),(99,99),(99,99)), 0,  6) -- 1251
,( 0, E,0,1,((16,19),(20,23),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 1252
,( 0, E,0,1,((18,21),(22,25),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 1253
,( 0, E,0,1,((20,23),(24,27),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 1254
,( 0, E,0,1,((22,25),(26,29),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 1255
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 1256
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 1257
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 1258
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 1259
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 1260
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 1261
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 1262
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 1263
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 1264
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 1265
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 1266
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 1267
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 1268
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 1269
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 1270
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 1271
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 1272
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 1273
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 1274
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 1275
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 1276
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 1277
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 1278
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 1279
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 1, 31) -- 1280
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 1, 31) -- 1281
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 1, 31) -- 1282
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 1, 31) -- 1283
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 1, 31) -- 1284
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 1, 31) -- 1285
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 1, 31) -- 1286
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 1, 31) -- 1287
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 1288
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 1289
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 1290
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 1291
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 1292
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 1293
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 1294
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 1295
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 31) -- 1296
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),(10,10)), 1, 31) -- 1297
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(11,11)), 1, 31) -- 1298
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(12,12)), 1, 31) -- 1299
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(13,13)), 1, 31) -- 1300
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(14,14)), 1, 31) -- 1301
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(15,15)), 1, 31) -- 1302
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(16,16)), 1, 31) -- 1303
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 31) -- 1304
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 31) -- 1305
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 1, 31) -- 1306
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 1, 31) -- 1307
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 1, 31) -- 1308
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 1, 31) -- 1309
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 1, 31) -- 1310
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 1, 31) -- 1311
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),(11,11)), 1, 31) -- 1312
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),(12,12)), 1, 31) -- 1313
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(13,13)), 1, 31) -- 1314
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(14,14)), 1, 31) -- 1315
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(15,15)), 1, 31) -- 1316
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(16,16)), 1, 31) -- 1317
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(17,17)), 1, 31) -- 1318
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(18,18)), 1, 31) -- 1319
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 31) -- 1320
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 31) -- 1321
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 31) -- 1322
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 31) -- 1323
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 31) -- 1324
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 31) -- 1325
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 31) -- 1326
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 31) -- 1327
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 30) -- 1328
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 30) -- 1329
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 30) -- 1330
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 30) -- 1331
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 30) -- 1332
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 30) -- 1333
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 30) -- 1334
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 30) -- 1335
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 30) -- 1336
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),(10,10)), 1, 30) -- 1337
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(11,11)), 1, 30) -- 1338
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(12,12)), 1, 30) -- 1339
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(13,13)), 1, 30) -- 1340
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(14,14)), 1, 30) -- 1341
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(15,15)), 1, 30) -- 1342
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(16,16)), 1, 30) -- 1343
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 30) -- 1344
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 30) -- 1345
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 30) -- 1346
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 30) -- 1347
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 30) -- 1348
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 30) -- 1349
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 30) -- 1350
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 30) -- 1351
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 29) -- 1352
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 29) -- 1353
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 29) -- 1354
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 29) -- 1355
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 29) -- 1356
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 29) -- 1357
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 29) -- 1358
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 29) -- 1359
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 28) -- 1360
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 28) -- 1361
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 28) -- 1362
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 28) -- 1363
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 28) -- 1364
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 28) -- 1365
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 28) -- 1366
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 28) -- 1367
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 28) -- 1368
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 28) -- 1369
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 28) -- 1370
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 28) -- 1371
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 28) -- 1372
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 28) -- 1373
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 28) -- 1374
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 28) -- 1375
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 1, 28) -- 1376
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 1, 28) -- 1377
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 1, 28) -- 1378
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 1, 28) -- 1379
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 1, 28) -- 1380
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 1, 28) -- 1381
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 1, 28) -- 1382
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 1, 28) -- 1383
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 27) -- 1384
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 27) -- 1385
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 27) -- 1386
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 27) -- 1387
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 27) -- 1388
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 27) -- 1389
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 27) -- 1390
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 27) -- 1391
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 26) -- 1392
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 26) -- 1393
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 26) -- 1394
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 26) -- 1395
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 26) -- 1396
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 26) -- 1397
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 26) -- 1398
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 26) -- 1399
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 25) -- 1400
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 25) -- 1401
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 25) -- 1402
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 25) -- 1403
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 25) -- 1404
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 25) -- 1405
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 25) -- 1406
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 25) -- 1407
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 24) -- 1408
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 24) -- 1409
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 24) -- 1410
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 24) -- 1411
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 24) -- 1412
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 24) -- 1413
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 24) -- 1414
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 24) -- 1415
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 1416
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 1417
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 1418
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 1419
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 1420
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 1421
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 1422
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 1423
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 22) -- 1424
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 22) -- 1425
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 22) -- 1426
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 22) -- 1427
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 22) -- 1428
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 22) -- 1429
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 22) -- 1430
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 22) -- 1431
,( 1, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 22) -- 1432
,( 1, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 22) -- 1433
,( 1, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 22) -- 1434
,( 1, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 22) -- 1435
,( 1, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 22) -- 1436
,( 1, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 22) -- 1437
,( 1, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 22) -- 1438
,( 1, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 22) -- 1439
,( 1, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 21) -- 1440
,( 1, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 21) -- 1441
,( 1, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 21) -- 1442
,( 1, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 21) -- 1443
,( 1, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 21) -- 1444
,( 1, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 21) -- 1445
,( 1, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 21) -- 1446
,( 1, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 21) -- 1447
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 21) -- 1448
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 21) -- 1449
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 21) -- 1450
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 21) -- 1451
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 21) -- 1452
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 21) -- 1453
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 21) -- 1454
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 21) -- 1455
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 1456
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 1457
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 1458
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 1459
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 1460
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 1461
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 1462
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 1463
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 20) -- 1464
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 20) -- 1465
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 20) -- 1466
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 20) -- 1467
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 20) -- 1468
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 20) -- 1469
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 20) -- 1470
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 20) -- 1471
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 20) -- 1472
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 20) -- 1473
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 20) -- 1474
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 20) -- 1475
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 20) -- 1476
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 20) -- 1477
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 20) -- 1478
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 20) -- 1479
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 1480
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 1481
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 1482
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 1483
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 1484
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 1485
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 1486
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 1487
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 19) -- 1488
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 19) -- 1489
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 19) -- 1490
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(19,19),(19,19),(10,10)), 1, 19) -- 1491
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(20,20),(20,20),(11,11)), 1, 19) -- 1492
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(21,21),(21,21),(12,12)), 1, 19) -- 1493
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(22,22),(22,22),(13,13)), 1, 19) -- 1494
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(23,23),(23,23),(14,14)), 1, 19) -- 1495
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 1496
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 1497
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 1498
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 1499
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 1500
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 1501
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 1502
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 1503
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 1504
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 1505
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 1506
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 1507
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 1508
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 1509
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 1510
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 1511
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 19) -- 1512
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 19) -- 1513
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 19) -- 1514
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 19) -- 1515
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 19) -- 1516
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 19) -- 1517
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 19) -- 1518
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 19) -- 1519
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 19) -- 1520
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 19) -- 1521
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(18,18),(18,18),(10,10)), 1, 19) -- 1522
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(19,19),(19,19),(11,11)), 1, 19) -- 1523
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(20,20),(20,20),(12,12)), 1, 19) -- 1524
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(21,21),(21,21),(13,13)), 1, 19) -- 1525
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(22,22),(22,22),(14,14)), 1, 19) -- 1526
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(23,23),(23,23),(15,15)), 1, 19) -- 1527
,( 1, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 19) -- 1528
,( 1, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 19) -- 1529
,( 1, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),(10,10)), 1, 19) -- 1530
,( 1, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(11,11)), 1, 19) -- 1531
,( 1, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(12,12)), 1, 19) -- 1532
,( 1, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(13,13)), 1, 19) -- 1533
,( 1, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(14,14)), 1, 19) -- 1534
,( 1, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(15,15)), 1, 19) -- 1535
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 1536
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 1537
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 1538
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 1539
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 1540
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 1541
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 1542
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 1543
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 1544
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 1545
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 1546
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 1547
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 1548
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 1549
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 1550
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 1551
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 1552
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 1553
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 1554
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 1555
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 1556
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 1557
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 1558
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 1559
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 18) -- 1560
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 18) -- 1561
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 18) -- 1562
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 18) -- 1563
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 18) -- 1564
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 18) -- 1565
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 18) -- 1566
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 18) -- 1567
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 18) -- 1568
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 18) -- 1569
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 18) -- 1570
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(19,19),(10,10)), 1, 18) -- 1571
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(20,20),(11,11)), 1, 18) -- 1572
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(21,21),(12,12)), 1, 18) -- 1573
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(22,22),(13,13)), 1, 18) -- 1574
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(23,23),(14,14)), 1, 18) -- 1575
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 17) -- 1576
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 17) -- 1577
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 17) -- 1578
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 17) -- 1579
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 17) -- 1580
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 17) -- 1581
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 17) -- 1582
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 17) -- 1583
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 1584
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 1585
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 1586
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 1587
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 1588
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 1589
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 1590
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 1591
,( 1, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 1592
,( 1, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 1593
,( 1, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 1594
,( 1, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 1595
,( 1, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 1596
,( 1, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 1597
,( 1, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 1598
,( 1, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 1599
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 1600
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 1601
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 1602
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 1603
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 1604
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 1605
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 1606
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 1607
,( 1, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 17) -- 1608
,( 1, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 17) -- 1609
,( 1, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 17) -- 1610
,( 1, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 17) -- 1611
,( 1, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 17) -- 1612
,( 1, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 17) -- 1613
,( 1, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 17) -- 1614
,( 1, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 17) -- 1615
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 16) -- 1616
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 16) -- 1617
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 16) -- 1618
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 16) -- 1619
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 16) -- 1620
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 16) -- 1621
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 16) -- 1622
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 16) -- 1623
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 16) -- 1624
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 16) -- 1625
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 16) -- 1626
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 16) -- 1627
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 16) -- 1628
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 16) -- 1629
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 16) -- 1630
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 16) -- 1631
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 16) -- 1632
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 16) -- 1633
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 16) -- 1634
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 16) -- 1635
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 16) -- 1636
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),(10,10)), 1, 16) -- 1637
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(11,11)), 1, 16) -- 1638
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(12,12)), 1, 16) -- 1639
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 1640
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 1641
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 1642
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 1643
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 1644
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 1645
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 1646
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 1647
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 1648
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 1649
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 1650
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 1651
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 1652
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 1653
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 1654
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 1655
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 1656
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 1657
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 1658
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 1659
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 1660
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 1661
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 1662
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 1663
,( 1, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 1664
,( 1, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 1665
,( 1, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 1666
,( 1, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 1667
,( 1, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 1668
,( 1, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 1669
,( 1, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 1670
,( 1, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 1671
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 15) -- 1672
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 15) -- 1673
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 15) -- 1674
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 15) -- 1675
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 15) -- 1676
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 15) -- 1677
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(10,10)), 1, 15) -- 1678
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(11,11)), 1, 15) -- 1679
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 1680
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 1681
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 1682
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 1683
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 1684
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 1685
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 1686
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 1687
,( 1, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 15) -- 1688
,( 1, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 15) -- 1689
,( 1, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),(10,10)), 1, 15) -- 1690
,( 1, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(11,11)), 1, 15) -- 1691
,( 1, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(12,12)), 1, 15) -- 1692
,( 1, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(13,13)), 1, 15) -- 1693
,( 1, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(14,14)), 1, 15) -- 1694
,( 1, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(15,15)), 1, 15) -- 1695
,( 1, E,0,0,((36,36),(27,27),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 1696
,( 1, E,0,0,((37,37),(28,28),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 1697
,( 1, E,0,0,((38,38),(29,29),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 1698
,( 1, E,0,0,((39,39),(30,30),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 1699
,( 1, E,0,0,((40,40),(31,31),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 1700
,( 1, E,0,0,((41,41),(32,32),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 1701
,( 1, E,0,0,((42,42),(33,33),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 1702
,( 1, E,0,0,((43,43),(34,34),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 1703
,( 1, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 1704
,( 1, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 1705
,( 1, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 1706
,( 1, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 1707
,( 1, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 1708
,( 1, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 1709
,( 1, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 1710
,( 1, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 1711
,( 1, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 1712
,( 1, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 1713
,( 1, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 1714
,( 1, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 1715
,( 1, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 1716
,( 1, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 1717
,( 1, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 1718
,( 1, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 1719
,( 1, E,0,0,((36,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 1720
,( 1, E,0,0,((38,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 1721
,( 1, E,0,0,((40,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 1722
,( 1, E,0,0,((42,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 1723
,( 1, E,0,0,((36,39),(28,29),( 1, 1),(15,15),(14,15),( 4, 7)), 1, 13) -- 1724
,( 1, E,0,0,((38,41),(30,31),( 3, 3),(17,17),(16,17),( 6, 9)), 1, 13) -- 1725
,( 1, E,0,0,((40,43),(32,33),( 5, 5),(19,19),(18,19),( 8,11)), 1, 13) -- 1726
,( 1, E,0,0,((42,45),(34,35),( 7, 7),(21,21),(20,21),(10,13)), 1, 13) -- 1727
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 1728
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 1729
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 1730
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 1731
,( 1, E,0,0,((38,38),(27,27),( 0, 0),(14,15),(12,13),( 2, 5)), 1, 12) -- 1732
,( 1, E,0,0,((40,40),(29,29),( 2, 2),(16,17),(14,15),( 4, 7)), 1, 12) -- 1733
,( 1, E,0,0,((42,42),(31,31),( 4, 4),(18,19),(16,17),( 6, 9)), 1, 12) -- 1734
,( 1, E,0,0,((44,44),(33,33),( 6, 6),(20,21),(18,19),( 8,11)), 1, 12) -- 1735
,( 1, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,13),( 2, 5)), 1, 12) -- 1736
,( 1, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,15),( 4, 7)), 1, 12) -- 1737
,( 1, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,17),( 6, 9)), 1, 12) -- 1738
,( 1, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,19),( 8,11)), 1, 12) -- 1739
,( 1, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 12) -- 1740
,( 1, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),( 8,11)), 1, 12) -- 1741
,( 1, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),(10,13)), 1, 12) -- 1742
,( 1, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(12,15)), 1, 12) -- 1743
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 1744
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 1745
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(10,13)), 1, 11) -- 1746
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(12,15)), 1, 11) -- 1747
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(12,13),(10,11),( 0, 3)), 1, 11) -- 1748
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(14,15),(12,13),( 2, 5)), 1, 11) -- 1749
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(16,17),(14,15),( 4, 7)), 1, 11) -- 1750
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(18,19),(16,17),( 6, 9)), 1, 11) -- 1751
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 1752
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 1753
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 1754
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 1755
,( 1, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),( 2, 5)), 1, 11) -- 1756
,( 1, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),( 4, 7)), 1, 11) -- 1757
,( 1, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),( 6, 9)), 1, 11) -- 1758
,( 1, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),( 8,11)), 1, 11) -- 1759
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(15,15),(14,14),( 4, 5)), 1, 11) -- 1760
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(17,17),(16,16),( 6, 7)), 1, 11) -- 1761
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(19,19),(18,18),( 8, 9)), 1, 11) -- 1762
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(21,21),(20,20),(10,11)), 1, 11) -- 1763
,( 1, E,0,0,((36,39),(26,27),( 0, 0),(14,14),(13,13),( 6, 9)), 1, 11) -- 1764
,( 1, E,0,0,((38,41),(28,29),( 2, 2),(16,16),(15,15),( 8,11)), 1, 11) -- 1765
,( 1, E,0,0,((40,43),(30,31),( 4, 4),(18,18),(17,17),(10,13)), 1, 11) -- 1766
,( 1, E,0,0,((42,45),(32,33),( 6, 6),(20,20),(19,19),(12,15)), 1, 11) -- 1767
,( 1, E,0,0,((40,43),(30,31),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 10) -- 1768
,( 1, E,0,0,((42,45),(32,33),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 10) -- 1769
,( 1, E,0,0,((44,47),(34,35),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 10) -- 1770
,( 1, E,0,0,((46,49),(36,37),( 7, 7),(20,21),(18,19),( 8,11)), 1, 10) -- 1771
,( 1, E,0,0,((40,43),(30,31),( 1, 1),(14,14),(11,11),( 0, 3)), 1, 10) -- 1772
,( 1, E,0,0,((42,45),(32,33),( 3, 3),(16,16),(13,13),( 2, 5)), 1, 10) -- 1773
,( 1, E,0,0,((44,47),(34,35),( 5, 5),(18,18),(15,15),( 4, 7)), 1, 10) -- 1774
,( 1, E,0,0,((46,49),(36,37),( 7, 7),(20,20),(17,17),( 6, 9)), 1, 10) -- 1775
,( 1, E,0,0,((38,41),(28,29),( 0, 0),(12,13),(10,11),( 4, 7)), 1, 10) -- 1776
,( 1, E,0,0,((40,43),(30,31),( 2, 2),(14,15),(12,13),( 6, 9)), 1, 10) -- 1777
,( 1, E,0,0,((42,45),(32,33),( 4, 4),(16,17),(14,15),( 8,11)), 1, 10) -- 1778
,( 1, E,0,0,((44,47),(34,35),( 6, 6),(18,19),(16,17),(10,13)), 1, 10) -- 1779
,( 1, E,0,0,((40,43),(30,30),( 0, 1),(13,13),(10,11),( 2, 5)), 1, 10) -- 1780
,( 1, E,0,0,((42,45),(32,32),( 2, 3),(15,15),(12,13),( 4, 7)), 1, 10) -- 1781
,( 1, E,0,0,((44,47),(34,34),( 4, 5),(17,17),(14,15),( 6, 9)), 1, 10) -- 1782
,( 1, E,0,0,((46,49),(36,36),( 6, 7),(19,19),(16,17),( 8,11)), 1, 10) -- 1783
,( 1, E,0,0,((40,43),(30,30),( 1, 1),(15,15),(14,14),( 6, 9)), 1, 10) -- 1784
,( 1, E,0,0,((42,45),(32,32),( 3, 3),(17,17),(16,16),( 8,11)), 1, 10) -- 1785
,( 1, E,0,0,((44,47),(34,34),( 5, 5),(19,19),(18,18),(10,13)), 1, 10) -- 1786
,( 1, E,0,0,((46,49),(36,36),( 7, 7),(21,21),(20,20),(12,15)), 1, 10) -- 1787
,( 1, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(11,11),( 0, 3)), 1, 10) -- 1788
,( 1, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(13,13),( 2, 5)), 1, 10) -- 1789
,( 1, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(15,15),( 4, 7)), 1, 10) -- 1790
,( 1, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(17,17),( 6, 9)), 1, 10) -- 1791
,( 1, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),( 6, 9)), 1, 10) -- 1792
,( 1, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),( 8,11)), 1, 10) -- 1793
,( 1, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),(10,13)), 1, 10) -- 1794
,( 1, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),(12,15)), 1, 10) -- 1795
,( 1, E,0,0,((40,43),(30,31),( 1, 1),(14,15),(12,13),( 6, 7)), 1, 10) -- 1796
,( 1, E,0,0,((42,45),(32,33),( 3, 3),(16,17),(14,15),( 8, 9)), 1, 10) -- 1797
,( 1, E,0,0,((44,47),(34,35),( 5, 5),(18,19),(16,17),(10,11)), 1, 10) -- 1798
,( 1, E,0,0,((46,49),(36,37),( 7, 7),(20,21),(18,19),(12,13)), 1, 10) -- 1799
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),( 8,11)), 1,  9) -- 1800
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(10,13)), 1,  9) -- 1801
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(12,15)), 1,  9) -- 1802
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(14,17)), 1,  9) -- 1803
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 1804
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 1805
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 1806
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 1807
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 1808
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 1809
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 1810
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 1811
,( 1, E,0,0,((40,43),(30,31),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 1812
,( 1, E,0,0,((42,45),(32,33),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 1813
,( 1, E,0,0,((44,47),(34,35),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 1814
,( 1, E,0,0,((46,49),(36,37),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 1815
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 8,11)), 1,  9) -- 1816
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(10,13)), 1,  9) -- 1817
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(12,15)), 1,  9) -- 1818
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(14,17)), 1,  9) -- 1819
,( 1, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(12,13),(10,13)), 1,  9) -- 1820
,( 1, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(14,15),(12,15)), 1,  9) -- 1821
,( 1, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(16,17),(14,17)), 1,  9) -- 1822
,( 1, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(18,19),(16,19)), 1,  9) -- 1823
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 0, 3)), 1,  9) -- 1824
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 2, 5)), 1,  9) -- 1825
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 4, 7)), 1,  9) -- 1826
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 6, 9)), 1,  9) -- 1827
,( 1, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 1828
,( 1, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 1829
,( 1, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 1830
,( 1, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 1831
,( 1, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 4, 7)), 1,  9) -- 1832
,( 1, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 6, 9)), 1,  9) -- 1833
,( 1, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 8,11)), 1,  9) -- 1834
,( 1, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),(10,13)), 1,  9) -- 1835
,( 1, E,0,0,((42,42),(29,29),( 0, 0),(12,13),(10,11),( 2, 5)), 1,  9) -- 1836
,( 1, E,0,0,((44,44),(31,31),( 2, 2),(14,15),(12,13),( 4, 7)), 1,  9) -- 1837
,( 1, E,0,0,((46,46),(33,33),( 4, 4),(16,17),(14,15),( 6, 9)), 1,  9) -- 1838
,( 1, E,0,0,((48,48),(35,35),( 6, 6),(18,19),(16,17),( 8,11)), 1,  9) -- 1839
,( 1, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(14,15),(14,17)), 1,  9) -- 1840
,( 1, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(16,17),(16,19)), 1,  9) -- 1841
,( 1, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(18,19),(18,21)), 1,  9) -- 1842
,( 1, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(20,21),(20,23)), 1,  9) -- 1843
,( 1, E,0,0,((40,43),(29,29),( 0, 1),(14,14),(12,13),(10,13)), 1,  9) -- 1844
,( 1, E,0,0,((42,45),(31,31),( 2, 3),(16,16),(14,15),(12,15)), 1,  9) -- 1845
,( 1, E,0,0,((44,47),(33,33),( 4, 5),(18,18),(16,17),(14,17)), 1,  9) -- 1846
,( 1, E,0,0,((46,49),(35,35),( 6, 7),(20,20),(18,19),(16,19)), 1,  9) -- 1847
,( 1, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(12,13),(12,15)), 1,  9) -- 1848
,( 1, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(14,15),(14,17)), 1,  9) -- 1849
,( 1, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(16,17),(16,19)), 1,  9) -- 1850
,( 1, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(18,19),(18,21)), 1,  9) -- 1851
,( 1, E,0,0,((42,42),(29,29),( 0, 0),(13,13),(12,13),( 6, 9)), 1,  9) -- 1852
,( 1, E,0,0,((44,44),(31,31),( 2, 2),(15,15),(14,15),( 8,11)), 1,  9) -- 1853
,( 1, E,0,0,((46,46),(33,33),( 4, 4),(17,17),(16,17),(10,13)), 1,  9) -- 1854
,( 1, E,0,0,((48,48),(35,35),( 6, 6),(19,19),(18,19),(12,15)), 1,  9) -- 1855
,( 1, E,0,0,((38,41),(28,29),( 0, 1),(13,13),(12,13),(14,17)), 1,  9) -- 1856
,( 1, E,0,0,((40,43),(30,31),( 2, 3),(15,15),(14,15),(16,19)), 1,  9) -- 1857
,( 1, E,0,0,((42,45),(32,33),( 4, 5),(17,17),(16,17),(18,21)), 1,  9) -- 1858
,( 1, E,0,0,((44,47),(34,35),( 6, 7),(19,19),(18,19),(20,23)), 1,  9) -- 1859
,( 1, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),(16,19)), 1,  9) -- 1860
,( 1, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),(18,21)), 1,  9) -- 1861
,( 1, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(20,23)), 1,  9) -- 1862
,( 1, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(22,23)), 1,  9) -- 1863
,( 1, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1,  9) -- 1864
,( 1, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 8,11)), 1,  9) -- 1865
,( 1, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(10,13)), 1,  9) -- 1866
,( 1, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(12,15)), 1,  9) -- 1867
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(13,13),(11,11),( 8,11)), 1,  9) -- 1868
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(15,15),(13,13),(10,13)), 1,  9) -- 1869
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(17,17),(15,15),(12,15)), 1,  9) -- 1870
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(19,19),(17,17),(14,17)), 1,  9) -- 1871
,( 1, E,0,0,((45,45),(32,32),( 1, 1),(13,13),(10,11),( 3, 3)), 1,  9) -- 1872
,( 1, E,0,0,((47,47),(34,34),( 3, 3),(15,15),(12,13),( 5, 5)), 1,  9) -- 1873
,( 1, E,0,0,((49,49),(36,36),( 5, 5),(17,17),(14,15),( 7, 7)), 1,  9) -- 1874
,( 1, E,0,0,((51,51),(38,38),( 7, 7),(19,19),(16,17),( 9, 9)), 1,  9) -- 1875
,( 1, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(12,13),( 6, 7)), 1,  9) -- 1876
,( 1, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(14,15),( 8, 9)), 1,  9) -- 1877
,( 1, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(16,17),(10,11)), 1,  9) -- 1878
,( 1, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(18,19),(12,13)), 1,  9) -- 1879
,( 1, E,0,0,((42,43),(30,30),( 0, 1),(13,13),(12,13),(12,15)), 1,  9) -- 1880
,( 1, E,0,0,((44,45),(32,32),( 2, 3),(15,15),(14,15),(14,17)), 1,  9) -- 1881
,( 1, E,0,0,((46,47),(34,34),( 4, 5),(17,17),(16,17),(16,19)), 1,  9) -- 1882
,( 1, E,0,0,((48,49),(36,36),( 6, 7),(19,19),(18,19),(18,21)), 1,  9) -- 1883
,( 1, E,0,0,((40,43),(30,30),( 0, 1),(13,13),(12,12),( 6, 9)), 1,  9) -- 1884
,( 1, E,0,0,((42,45),(32,32),( 2, 3),(15,15),(14,14),( 8,11)), 1,  9) -- 1885
,( 1, E,0,0,((44,47),(34,34),( 4, 5),(17,17),(16,16),(10,13)), 1,  9) -- 1886
,( 1, E,0,0,((46,49),(36,36),( 6, 7),(19,19),(18,18),(12,15)), 1,  9) -- 1887
,( 1, E,0,0,((40,43),(29,29),( 0, 0),(12,12),( 8, 9),( 0, 3)), 1,  9) -- 1888
,( 1, E,0,0,((42,45),(31,31),( 2, 2),(14,14),(10,11),( 2, 5)), 1,  9) -- 1889
,( 1, E,0,0,((44,47),(33,33),( 4, 4),(16,16),(12,13),( 4, 7)), 1,  9) -- 1890
,( 1, E,0,0,((46,49),(35,35),( 6, 6),(18,18),(14,15),( 6, 9)), 1,  9) -- 1891
,( 1, E,0,0,((38,41),(28,29),( 0, 0),(14,14),(12,13),(14,17)), 1,  9) -- 1892
,( 1, E,0,0,((40,43),(30,31),( 2, 2),(16,16),(14,15),(16,19)), 1,  9) -- 1893
,( 1, E,0,0,((42,45),(32,33),( 4, 4),(18,18),(16,17),(18,21)), 1,  9) -- 1894
,( 1, E,0,0,((44,47),(34,35),( 6, 6),(20,20),(18,19),(20,23)), 1,  9) -- 1895
,( 1, E,0,0,((42,45),(31,31),( 1, 1),(14,14),(10,11),( 0, 3)), 1,  9) -- 1896
,( 1, E,0,0,((44,47),(33,33),( 3, 3),(16,16),(12,13),( 2, 5)), 1,  9) -- 1897
,( 1, E,0,0,((46,49),(35,35),( 5, 5),(18,18),(14,15),( 4, 7)), 1,  9) -- 1898
,( 1, E,0,0,((48,51),(37,37),( 7, 7),(20,20),(16,17),( 6, 9)), 1,  9) -- 1899
,( 1, E,0,0,((40,43),(29,29),( 0, 0),(12,13),(11,11),(10,10)), 1,  9) -- 1900
,( 1, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(13,13),(12,12)), 1,  9) -- 1901
,( 1, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(15,15),(14,14)), 1,  9) -- 1902
,( 1, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(17,17),(16,16)), 1,  9) -- 1903
,( 1, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(10,13),(16,19)), 1,  8) -- 1904
,( 1, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(12,15),(18,21)), 1,  8) -- 1905
,( 1, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(14,17),(20,23)), 1,  8) -- 1906
,( 1, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(16,19),(22,23)), 1,  8) -- 1907
,( 1, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(16,16)), 1,  8) -- 1908
,( 1, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(18,18)), 1,  8) -- 1909
,( 1, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(20,20)), 1,  8) -- 1910
,( 1, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(22,22)), 1,  8) -- 1911
,( 1, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 6, 9),( 0, 3)), 1,  8) -- 1912
,( 1, E,0,0,((46,49),(32,35),( 2, 3),(12,15),( 8,11),( 2, 5)), 1,  8) -- 1913
,( 1, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(10,13),( 4, 7)), 1,  8) -- 1914
,( 1, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(12,15),( 6, 9)), 1,  8) -- 1915
,( 1, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(12,15),(99,99)), 1,  8) -- 1916
,( 1, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(14,17),(99,99)), 1,  8) -- 1917
,( 1, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(16,19),(99,99)), 1,  8) -- 1918
,( 1, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(18,21),(99,99)), 1,  8) -- 1919
,( 1, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(16,19),(99,99)), 1,  7) -- 1920
,( 1, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(18,21),(99,99)), 1,  7) -- 1921
,( 1, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(20,23),(99,99)), 1,  7) -- 1922
,( 1, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(22,25),(99,99)), 1,  7) -- 1923
,( 1, E,0,0,((48,51),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 1924
,( 1, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 1925
,( 1, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 1926
,( 1, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 1927
,( 1, E,0,1,((48,51),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 1928
,( 1, E,0,1,((50,53),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 1929
,( 1, E,0,1,((52,55),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 1930
,( 1, E,0,1,((54,57),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 1931
,( 1, E,0,1,((46,49),(30,33),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 1932
,( 1, E,0,1,((48,51),(32,35),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 1933
,( 1, E,0,1,((50,53),(34,37),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 1934
,( 1, E,0,1,((52,55),(36,39),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 1935
,( 1, E,0,1,((50,53),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  6) -- 1936
,( 1, E,0,1,((52,55),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  6) -- 1937
,( 1, E,0,1,((54,57),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  6) -- 1938
,( 1, E,0,1,((56,59),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  6) -- 1939
,( 1, E,0,1,((38,41),(24,27),( 0, 1),(18,21),(99,99),(99,99)), 1,  5) -- 1940
,( 1, E,0,1,((40,43),(26,29),( 2, 3),(20,23),(99,99),(99,99)), 1,  5) -- 1941
,( 1, E,0,1,((42,45),(28,31),( 4, 5),(22,25),(99,99),(99,99)), 1,  5) -- 1942
,( 1, E,0,1,((44,47),(30,33),( 6, 7),(24,27),(99,99),(99,99)), 1,  5) -- 1943
,( 1, E,0,1,((46,49),(30,33),( 0, 1),(20,23),(99,99),(99,99)), 1,  5) -- 1944
,( 1, E,0,1,((48,51),(32,35),( 2, 3),(22,25),(99,99),(99,99)), 1,  5) -- 1945
,( 1, E,0,1,((50,53),(34,37),( 4, 5),(24,27),(99,99),(99,99)), 1,  5) -- 1946
,( 1, E,0,1,((52,55),(36,39),( 6, 7),(26,29),(99,99),(99,99)), 1,  5) -- 1947
,( 1, E,0,1,((40,43),(28,28),( 1, 1),(20,21),(99,99),(99,99)), 1,  5) -- 1948
,( 1, E,0,1,((42,45),(30,30),( 3, 3),(22,23),(99,99),(99,99)), 1,  5) -- 1949
,( 1, E,0,1,((44,47),(32,32),( 5, 5),(24,25),(99,99),(99,99)), 1,  5) -- 1950
,( 1, E,0,1,((46,49),(34,34),( 7, 7),(26,27),(99,99),(99,99)), 1,  5) -- 1951
,( 1, E,0,1,((26,29),(20,21),( 0, 1),(24,27),(99,99),(99,99)), 1,  5) -- 1952
,( 1, E,0,1,((28,31),(22,23),( 2, 3),(26,29),(99,99),(99,99)), 1,  5) -- 1953
,( 1, E,0,1,((30,33),(24,25),( 4, 5),(28,31),(99,99),(99,99)), 1,  5) -- 1954
,( 1, E,0,1,((32,35),(26,27),( 6, 7),(30,33),(99,99),(99,99)), 1,  5) -- 1955
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 1956
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 1957
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 1958
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 1959
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 1960
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 1961
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 1962
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 1963
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 1964
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 1965
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 1966
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 1967
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 1968
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 1969
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 1970
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 1971
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 1972
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 1973
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 1974
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 1975
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 1976
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 1977
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 1978
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 1979
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 1980
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 1981
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 1982
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 1983
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 1984
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 1985
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 1986
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 1987
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 1988
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 1989
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 1990
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 1991
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 1992
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 1993
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 1994
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 1995
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 1996
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 1997
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 1998
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 1999
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 2000
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 2001
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 2002
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 2003
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 31) -- 2004
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),(10,10)), 0, 31) -- 2005
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(11,11)), 0, 31) -- 2006
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(12,12)), 0, 31) -- 2007
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(13,13)), 0, 31) -- 2008
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(14,14)), 0, 31) -- 2009
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(15,15)), 0, 31) -- 2010
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(16,16)), 0, 31) -- 2011
,( 1, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 2012
,( 1, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 2013
,( 1, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 2014
,( 1, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 2015
,( 1, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 2016
,( 1, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 2017
,( 1, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 2018
,( 1, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 2019
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 2020
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 2021
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 2022
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 2023
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 2024
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 2025
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 2026
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 2027
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 2028
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 2029
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 2030
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 2031
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 2032
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 2033
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 2034
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 2035
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 30) -- 2036
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 30) -- 2037
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 30) -- 2038
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 30) -- 2039
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 30) -- 2040
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 30) -- 2041
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 30) -- 2042
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 30) -- 2043
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 30) -- 2044
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 30) -- 2045
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 30) -- 2046
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 30) -- 2047
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 30) -- 2048
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 30) -- 2049
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 30) -- 2050
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 30) -- 2051
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 28) -- 2052
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 28) -- 2053
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 28) -- 2054
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 28) -- 2055
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 28) -- 2056
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 28) -- 2057
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 28) -- 2058
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 28) -- 2059
,( 1, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 27) -- 2060
,( 1, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 27) -- 2061
,( 1, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 27) -- 2062
,( 1, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 27) -- 2063
,( 1, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 27) -- 2064
,( 1, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 27) -- 2065
,( 1, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 27) -- 2066
,( 1, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 27) -- 2067
,( 1, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 26) -- 2068
,( 1, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 26) -- 2069
,( 1, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 26) -- 2070
,( 1, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 26) -- 2071
,( 1, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 26) -- 2072
,( 1, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 26) -- 2073
,( 1, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 26) -- 2074
,( 1, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 26) -- 2075
,( 1, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 26) -- 2076
,( 1, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 26) -- 2077
,( 1, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 26) -- 2078
,( 1, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 26) -- 2079
,( 1, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 26) -- 2080
,( 1, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 26) -- 2081
,( 1, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 26) -- 2082
,( 1, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 26) -- 2083
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 25) -- 2084
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 25) -- 2085
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 25) -- 2086
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 25) -- 2087
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 25) -- 2088
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 25) -- 2089
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 25) -- 2090
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 25) -- 2091
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(13,13)), 0, 24) -- 2092
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(14,14)), 0, 24) -- 2093
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(15,15)), 0, 24) -- 2094
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(16,16)), 0, 24) -- 2095
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(17,17)), 0, 24) -- 2096
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(18,18)), 0, 24) -- 2097
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(19,19)), 0, 24) -- 2098
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(20,20)), 0, 24) -- 2099
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(17,17),( 9, 9)), 0, 24) -- 2100
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(18,18),(10,10)), 0, 24) -- 2101
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(19,19),(11,11)), 0, 24) -- 2102
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(20,20),(12,12)), 0, 24) -- 2103
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(21,21),(13,13)), 0, 24) -- 2104
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(22,22),(14,14)), 0, 24) -- 2105
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(23,23),(15,15)), 0, 24) -- 2106
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(24,24),(16,16)), 0, 24) -- 2107
,( 1, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 24) -- 2108
,( 1, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 24) -- 2109
,( 1, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 24) -- 2110
,( 1, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 24) -- 2111
,( 1, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 24) -- 2112
,( 1, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 24) -- 2113
,( 1, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 24) -- 2114
,( 1, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 24) -- 2115
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 23) -- 2116
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 23) -- 2117
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 23) -- 2118
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 23) -- 2119
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 23) -- 2120
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 23) -- 2121
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 23) -- 2122
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 23) -- 2123
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 23) -- 2124
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 23) -- 2125
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 23) -- 2126
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 23) -- 2127
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 23) -- 2128
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 23) -- 2129
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 23) -- 2130
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 23) -- 2131
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 23) -- 2132
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 23) -- 2133
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 23) -- 2134
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 23) -- 2135
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 23) -- 2136
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 23) -- 2137
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 23) -- 2138
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 23) -- 2139
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 22) -- 2140
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 22) -- 2141
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 22) -- 2142
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 22) -- 2143
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 22) -- 2144
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 22) -- 2145
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 22) -- 2146
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 22) -- 2147
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 21) -- 2148
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 21) -- 2149
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 21) -- 2150
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 21) -- 2151
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 21) -- 2152
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 21) -- 2153
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 21) -- 2154
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 21) -- 2155
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 2156
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 2157
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 2158
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 2159
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 2160
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 2161
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 2162
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 2163
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 20) -- 2164
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 20) -- 2165
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 20) -- 2166
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 20) -- 2167
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 20) -- 2168
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 20) -- 2169
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 20) -- 2170
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 20) -- 2171
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 2172
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 2173
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 2174
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 2175
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 2176
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 2177
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 2178
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 2179
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 2180
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 2181
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 2182
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 2183
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 2184
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 2185
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 2186
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 2187
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 20) -- 2188
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(10,10)), 0, 20) -- 2189
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(11,11)), 0, 20) -- 2190
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(12,12)), 0, 20) -- 2191
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(13,13)), 0, 20) -- 2192
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(14,14)), 0, 20) -- 2193
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(15,15)), 0, 20) -- 2194
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(16,16)), 0, 20) -- 2195
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(11,11)), 0, 19) -- 2196
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(12,12)), 0, 19) -- 2197
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(13,13)), 0, 19) -- 2198
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(14,14)), 0, 19) -- 2199
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(15,15)), 0, 19) -- 2200
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(16,16)), 0, 19) -- 2201
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(17,17)), 0, 19) -- 2202
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(18,18)), 0, 19) -- 2203
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),(11,11)), 0, 19) -- 2204
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(12,12)), 0, 19) -- 2205
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(13,13)), 0, 19) -- 2206
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(14,14)), 0, 19) -- 2207
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(15,15)), 0, 19) -- 2208
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(16,16)), 0, 19) -- 2209
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(17,17)), 0, 19) -- 2210
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(18,18)), 0, 19) -- 2211
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 2212
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 2213
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 2214
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 2215
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 2216
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 2217
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 2218
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 2219
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 19) -- 2220
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 19) -- 2221
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 19) -- 2222
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 19) -- 2223
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 19) -- 2224
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 19) -- 2225
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 19) -- 2226
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 19) -- 2227
,( 1, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(18,18),(11,11)), 0, 19) -- 2228
,( 1, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(19,19),(12,12)), 0, 19) -- 2229
,( 1, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(20,20),(13,13)), 0, 19) -- 2230
,( 1, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(21,21),(14,14)), 0, 19) -- 2231
,( 1, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(22,22),(15,15)), 0, 19) -- 2232
,( 1, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(23,23),(16,16)), 0, 19) -- 2233
,( 1, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(24,24),(17,17)), 0, 19) -- 2234
,( 1, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(25,25),(18,18)), 0, 19) -- 2235
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),(13,13)), 0, 19) -- 2236
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(14,14)), 0, 19) -- 2237
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(15,15)), 0, 19) -- 2238
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(16,16)), 0, 19) -- 2239
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(17,17)), 0, 19) -- 2240
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(18,18)), 0, 19) -- 2241
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(19,19)), 0, 19) -- 2242
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(20,20)), 0, 19) -- 2243
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 2244
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 2245
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 2246
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 2247
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 2248
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 2249
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 2250
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 2251
,( 1, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 19) -- 2252
,( 1, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(10,10)), 0, 19) -- 2253
,( 1, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(11,11)), 0, 19) -- 2254
,( 1, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(12,12)), 0, 19) -- 2255
,( 1, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(13,13)), 0, 19) -- 2256
,( 1, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(14,14)), 0, 19) -- 2257
,( 1, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(15,15)), 0, 19) -- 2258
,( 1, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(16,16)), 0, 19) -- 2259
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 2260
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 2261
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 2262
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 2263
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 2264
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 2265
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 2266
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 2267
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 2268
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 2269
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 2270
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 2271
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 2272
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 2273
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 2274
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 2275
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 18) -- 2276
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 18) -- 2277
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 18) -- 2278
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 18) -- 2279
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 18) -- 2280
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 18) -- 2281
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 18) -- 2282
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 18) -- 2283
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 18) -- 2284
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 18) -- 2285
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 18) -- 2286
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 18) -- 2287
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 18) -- 2288
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 18) -- 2289
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 18) -- 2290
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 18) -- 2291
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 2292
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 2293
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 2294
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 2295
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 2296
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 2297
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 2298
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 2299
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 18) -- 2300
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 18) -- 2301
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 18) -- 2302
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 18) -- 2303
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 18) -- 2304
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 18) -- 2305
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 18) -- 2306
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 18) -- 2307
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(13,13)), 0, 18) -- 2308
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(14,14)), 0, 18) -- 2309
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(15,15)), 0, 18) -- 2310
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(16,16)), 0, 18) -- 2311
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(17,17)), 0, 18) -- 2312
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(18,18)), 0, 18) -- 2313
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(19,19)), 0, 18) -- 2314
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(20,20)), 0, 18) -- 2315
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 18) -- 2316
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 18) -- 2317
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 18) -- 2318
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 18) -- 2319
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 18) -- 2320
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 18) -- 2321
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 18) -- 2322
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 18) -- 2323
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 2324
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 2325
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 2326
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 2327
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 2328
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 2329
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 2330
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 2331
,( 1, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 17) -- 2332
,( 1, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 17) -- 2333
,( 1, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 17) -- 2334
,( 1, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 17) -- 2335
,( 1, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 17) -- 2336
,( 1, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 17) -- 2337
,( 1, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 17) -- 2338
,( 1, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 17) -- 2339
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 17) -- 2340
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 17) -- 2341
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 17) -- 2342
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 17) -- 2343
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 17) -- 2344
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 17) -- 2345
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 17) -- 2346
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 17) -- 2347
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 17) -- 2348
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 17) -- 2349
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 17) -- 2350
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 17) -- 2351
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 17) -- 2352
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 17) -- 2353
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 17) -- 2354
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 17) -- 2355
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 2356
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 2357
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 2358
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 2359
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 2360
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 2361
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 2362
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 2363
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 17) -- 2364
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 17) -- 2365
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 17) -- 2366
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 17) -- 2367
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 17) -- 2368
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 17) -- 2369
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 17) -- 2370
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 17) -- 2371
,( 1, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 2372
,( 1, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 2373
,( 1, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 2374
,( 1, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 2375
,( 1, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 2376
,( 1, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 2377
,( 1, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 2378
,( 1, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 2379
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(14,14)), 0, 17) -- 2380
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(15,15)), 0, 17) -- 2381
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(16,16)), 0, 17) -- 2382
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(17,17)), 0, 17) -- 2383
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(18,18)), 0, 17) -- 2384
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(19,19)), 0, 17) -- 2385
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(20,20)), 0, 17) -- 2386
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(21,21)), 0, 17) -- 2387
,( 1, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 17) -- 2388
,( 1, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 17) -- 2389
,( 1, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 17) -- 2390
,( 1, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 17) -- 2391
,( 1, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 17) -- 2392
,( 1, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 17) -- 2393
,( 1, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 17) -- 2394
,( 1, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 17) -- 2395
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(14,14)), 0, 17) -- 2396
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(15,15)), 0, 17) -- 2397
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(16,16)), 0, 17) -- 2398
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(17,17)), 0, 17) -- 2399
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(18,18)), 0, 17) -- 2400
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(19,19)), 0, 17) -- 2401
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(20,20)), 0, 17) -- 2402
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(21,21)), 0, 17) -- 2403
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 2404
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 2405
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 2406
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 2407
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 2408
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 2409
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 2410
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 2411
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 2412
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 2413
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 2414
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 2415
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 2416
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 2417
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 2418
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 2419
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 2420
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 2421
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 2422
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 2423
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 2424
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 2425
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 2426
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 2427
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(12,12)), 0, 16) -- 2428
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(13,13)), 0, 16) -- 2429
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(14,14)), 0, 16) -- 2430
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(15,15)), 0, 16) -- 2431
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(16,16)), 0, 16) -- 2432
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(17,17)), 0, 16) -- 2433
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(18,18)), 0, 16) -- 2434
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(19,19)), 0, 16) -- 2435
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(12,12)), 0, 16) -- 2436
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(13,13)), 0, 16) -- 2437
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(14,14)), 0, 16) -- 2438
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(15,15)), 0, 16) -- 2439
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(16,16)), 0, 16) -- 2440
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(17,17)), 0, 16) -- 2441
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(18,18)), 0, 16) -- 2442
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(19,19)), 0, 16) -- 2443
,( 1, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 16) -- 2444
,( 1, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 16) -- 2445
,( 1, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 16) -- 2446
,( 1, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 16) -- 2447
,( 1, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 16) -- 2448
,( 1, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 16) -- 2449
,( 1, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 16) -- 2450
,( 1, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 16) -- 2451
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(13,13)), 0, 16) -- 2452
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(14,14)), 0, 16) -- 2453
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(15,15)), 0, 16) -- 2454
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(16,16)), 0, 16) -- 2455
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(17,17)), 0, 16) -- 2456
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(18,18)), 0, 16) -- 2457
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(19,19)), 0, 16) -- 2458
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(20,20)), 0, 16) -- 2459
,( 1, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 16) -- 2460
,( 1, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(10,10)), 0, 16) -- 2461
,( 1, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(11,11)), 0, 16) -- 2462
,( 1, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(12,12)), 0, 16) -- 2463
,( 1, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(13,13)), 0, 16) -- 2464
,( 1, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(14,14)), 0, 16) -- 2465
,( 1, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(15,15)), 0, 16) -- 2466
,( 1, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(16,16)), 0, 16) -- 2467
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 2468
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 2469
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 2470
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 2471
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 2472
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 2473
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 2474
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 2475
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(19,19),(11,11)), 0, 15) -- 2476
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(20,20),(12,12)), 0, 15) -- 2477
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(21,21),(13,13)), 0, 15) -- 2478
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(22,22),(14,14)), 0, 15) -- 2479
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(23,23),(15,15)), 0, 15) -- 2480
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(24,24),(16,16)), 0, 15) -- 2481
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(25,25),(17,17)), 0, 15) -- 2482
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(26,26),(18,18)), 0, 15) -- 2483
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(13,13)), 0, 15) -- 2484
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(14,14)), 0, 15) -- 2485
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(15,15)), 0, 15) -- 2486
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(16,16)), 0, 15) -- 2487
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(17,17)), 0, 15) -- 2488
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(18,18)), 0, 15) -- 2489
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(19,19)), 0, 15) -- 2490
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(20,20)), 0, 15) -- 2491
,( 1, E,0,0,((28,28),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 2492
,( 1, E,0,0,((29,29),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 2493
,( 1, E,0,0,((30,30),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 2494
,( 1, E,0,0,((31,31),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 2495
,( 1, E,0,0,((32,32),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 2496
,( 1, E,0,0,((33,33),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 2497
,( 1, E,0,0,((34,34),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 2498
,( 1, E,0,0,((35,35),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 2499
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(12,12)), 0, 15) -- 2500
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(13,13)), 0, 15) -- 2501
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(14,14)), 0, 15) -- 2502
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(15,15)), 0, 15) -- 2503
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(16,16)), 0, 15) -- 2504
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(17,17)), 0, 15) -- 2505
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(18,18)), 0, 15) -- 2506
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(19,19)), 0, 15) -- 2507
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(13,13)), 0, 15) -- 2508
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(14,14)), 0, 15) -- 2509
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(15,15)), 0, 15) -- 2510
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(16,16)), 0, 15) -- 2511
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(17,17)), 0, 15) -- 2512
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(18,18)), 0, 15) -- 2513
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(19,19)), 0, 15) -- 2514
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(20,20)), 0, 15) -- 2515
,( 1, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(10,10)), 0, 15) -- 2516
,( 1, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(11,11)), 0, 15) -- 2517
,( 1, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(12,12)), 0, 15) -- 2518
,( 1, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(13,13)), 0, 15) -- 2519
,( 1, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(14,14)), 0, 15) -- 2520
,( 1, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(15,15)), 0, 15) -- 2521
,( 1, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(16,16)), 0, 15) -- 2522
,( 1, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(17,17)), 0, 15) -- 2523
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 2524
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 2525
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 2526
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 2527
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 2528
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 2529
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 2530
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 2531
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(14,14)), 0, 15) -- 2532
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(15,15)), 0, 15) -- 2533
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(16,16)), 0, 15) -- 2534
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(17,17)), 0, 15) -- 2535
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(18,18)), 0, 15) -- 2536
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(19,19)), 0, 15) -- 2537
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(20,20)), 0, 15) -- 2538
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(21,21)), 0, 15) -- 2539
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 15) -- 2540
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 15) -- 2541
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 15) -- 2542
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 15) -- 2543
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 15) -- 2544
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 15) -- 2545
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 15) -- 2546
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 15) -- 2547
,( 1, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(19,19),(12,12)), 0, 15) -- 2548
,( 1, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(20,20),(13,13)), 0, 15) -- 2549
,( 1, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(21,21),(14,14)), 0, 15) -- 2550
,( 1, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(22,22),(15,15)), 0, 15) -- 2551
,( 1, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(23,23),(16,16)), 0, 15) -- 2552
,( 1, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(24,24),(17,17)), 0, 15) -- 2553
,( 1, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(25,25),(18,18)), 0, 15) -- 2554
,( 1, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(26,26),(19,19)), 0, 15) -- 2555
,( 1, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 2556
,( 1, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 2557
,( 1, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 2558
,( 1, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 2559
,( 1, E,0,0,((26,29),(22,23),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 2560
,( 1, E,0,0,((28,31),(24,25),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 2561
,( 1, E,0,0,((30,33),(26,27),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 2562
,( 1, E,0,0,((32,35),(28,29),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 2563
,( 1, E,0,0,((28,31),(24,24),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 2564
,( 1, E,0,0,((30,33),(26,26),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 2565
,( 1, E,0,0,((32,35),(28,28),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 2566
,( 1, E,0,0,((34,37),(30,30),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 2567
,( 1, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(20,20),(12,15)), 0, 14) -- 2568
,( 1, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(22,22),(14,17)), 0, 14) -- 2569
,( 1, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(24,24),(16,19)), 0, 14) -- 2570
,( 1, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(26,26),(18,21)), 0, 14) -- 2571
,( 1, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(14,17)), 0, 14) -- 2572
,( 1, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(16,19)), 0, 14) -- 2573
,( 1, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(18,21)), 0, 14) -- 2574
,( 1, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(20,23)), 0, 14) -- 2575
,( 1, E,0,0,((26,27),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 13) -- 2576
,( 1, E,0,0,((28,29),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 13) -- 2577
,( 1, E,0,0,((30,31),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 13) -- 2578
,( 1, E,0,0,((32,33),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 13) -- 2579
,( 1, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(14,17)), 0, 13) -- 2580
,( 1, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(16,19)), 0, 13) -- 2581
,( 1, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(18,21)), 0, 13) -- 2582
,( 1, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(20,23)), 0, 13) -- 2583
,( 1, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(10,13)), 0, 13) -- 2584
,( 1, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(12,15)), 0, 13) -- 2585
,( 1, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(14,17)), 0, 13) -- 2586
,( 1, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(16,19)), 0, 13) -- 2587
,( 1, E,0,0,((28,29),(22,23),( 1, 1),(18,18),(19,19),(10,13)), 0, 13) -- 2588
,( 1, E,0,0,((30,31),(24,25),( 3, 3),(20,20),(21,21),(12,15)), 0, 13) -- 2589
,( 1, E,0,0,((32,33),(26,27),( 5, 5),(22,22),(23,23),(14,17)), 0, 13) -- 2590
,( 1, E,0,0,((34,35),(28,29),( 7, 7),(24,24),(25,25),(16,19)), 0, 13) -- 2591
,( 1, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(12,15)), 0, 12) -- 2592
,( 1, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(14,17)), 0, 12) -- 2593
,( 1, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(16,19)), 0, 12) -- 2594
,( 1, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(18,21)), 0, 12) -- 2595
,( 1, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 2596
,( 1, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 2597
,( 1, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 2598
,( 1, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 2599
,( 1, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(22,23),(14,17)), 0, 12) -- 2600
,( 1, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(24,25),(16,19)), 0, 12) -- 2601
,( 1, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(26,27),(18,21)), 0, 12) -- 2602
,( 1, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(28,29),(20,23)), 0, 12) -- 2603
,( 1, E,0,0,((24,27),(21,21),( 0, 0),(16,17),(18,19),( 8,11)), 0, 12) -- 2604
,( 1, E,0,0,((26,29),(23,23),( 2, 2),(18,19),(20,21),(10,13)), 0, 12) -- 2605
,( 1, E,0,0,((28,31),(25,25),( 4, 4),(20,21),(22,23),(12,15)), 0, 12) -- 2606
,( 1, E,0,0,((30,33),(27,27),( 6, 6),(22,23),(24,25),(14,17)), 0, 12) -- 2607
,( 1, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 12) -- 2608
,( 1, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 12) -- 2609
,( 1, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 12) -- 2610
,( 1, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 12) -- 2611
,( 1, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 2612
,( 1, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 2613
,( 1, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 2614
,( 1, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 2615
,( 1, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(20,21),(10,13)), 0, 11) -- 2616
,( 1, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(22,23),(12,15)), 0, 11) -- 2617
,( 1, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(24,25),(14,17)), 0, 11) -- 2618
,( 1, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(26,27),(16,19)), 0, 11) -- 2619
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(12,15)), 0, 11) -- 2620
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(14,17)), 0, 11) -- 2621
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(16,19)), 0, 11) -- 2622
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(18,21)), 0, 11) -- 2623
,( 1, E,0,0,((24,27),(22,23),( 1, 1),(19,19),(22,23),(12,15)), 0, 11) -- 2624
,( 1, E,0,0,((26,29),(24,25),( 3, 3),(21,21),(24,25),(14,17)), 0, 11) -- 2625
,( 1, E,0,0,((28,31),(26,27),( 5, 5),(23,23),(26,27),(16,19)), 0, 11) -- 2626
,( 1, E,0,0,((30,33),(28,29),( 7, 7),(25,25),(28,29),(18,21)), 0, 11) -- 2627
,( 1, E,0,0,((24,25),(20,21),( 0, 0),(17,17),(19,19),(10,13)), 0, 11) -- 2628
,( 1, E,0,0,((26,27),(22,23),( 2, 2),(19,19),(21,21),(12,15)), 0, 11) -- 2629
,( 1, E,0,0,((28,29),(24,25),( 4, 4),(21,21),(23,23),(14,17)), 0, 11) -- 2630
,( 1, E,0,0,((30,31),(26,27),( 6, 6),(23,23),(25,25),(16,19)), 0, 11) -- 2631
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(16,19)), 0, 11) -- 2632
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(18,21)), 0, 11) -- 2633
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(20,23)), 0, 11) -- 2634
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(22,23)), 0, 11) -- 2635
,( 1, E,0,0,((24,27),(22,23),( 1, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 2636
,( 1, E,0,0,((26,29),(24,25),( 3, 3),(20,21),(22,23),(10,13)), 0, 11) -- 2637
,( 1, E,0,0,((28,31),(26,27),( 5, 5),(22,23),(24,25),(12,15)), 0, 11) -- 2638
,( 1, E,0,0,((30,33),(28,29),( 7, 7),(24,25),(26,27),(14,17)), 0, 11) -- 2639
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,18),(20,21),(16,19)), 0, 11) -- 2640
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,20),(22,23),(18,21)), 0, 11) -- 2641
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,22),(24,25),(20,23)), 0, 11) -- 2642
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,24),(26,27),(22,23)), 0, 11) -- 2643
,( 1, E,0,0,((24,27),(22,23),( 1, 1),(19,19),(22,23),(16,19)), 0, 11) -- 2644
,( 1, E,0,0,((26,29),(24,25),( 3, 3),(21,21),(24,25),(18,21)), 0, 11) -- 2645
,( 1, E,0,0,((28,31),(26,27),( 5, 5),(23,23),(26,27),(20,23)), 0, 11) -- 2646
,( 1, E,0,0,((30,33),(28,29),( 7, 7),(25,25),(28,29),(22,23)), 0, 11) -- 2647
,( 1, E,0,0,((23,23),(20,20),( 0, 0),(18,18),(20,21),(10,13)), 0, 11) -- 2648
,( 1, E,0,0,((25,25),(22,22),( 2, 2),(20,20),(22,23),(12,15)), 0, 11) -- 2649
,( 1, E,0,0,((27,27),(24,24),( 4, 4),(22,22),(24,25),(14,17)), 0, 11) -- 2650
,( 1, E,0,0,((29,29),(26,26),( 6, 6),(24,24),(26,27),(16,19)), 0, 11) -- 2651
,( 1, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 2652
,( 1, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 2653
,( 1, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 2654
,( 1, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 2655
,( 1, E,0,0,((20,23),(19,19),( 0, 1),(18,19),(20,21),(10,13)), 0, 10) -- 2656
,( 1, E,0,0,((22,25),(21,21),( 2, 3),(20,21),(22,23),(12,15)), 0, 10) -- 2657
,( 1, E,0,0,((24,27),(23,23),( 4, 5),(22,23),(24,25),(14,17)), 0, 10) -- 2658
,( 1, E,0,0,((26,29),(25,25),( 6, 7),(24,25),(26,27),(16,19)), 0, 10) -- 2659
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 2660
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 2661
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 2662
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 2663
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(17,17),(18,19),( 6, 9)), 0, 10) -- 2664
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(19,19),(20,21),( 8,11)), 0, 10) -- 2665
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(21,21),(22,23),(10,13)), 0, 10) -- 2666
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(23,23),(24,25),(12,15)), 0, 10) -- 2667
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),( 8,11)), 0, 10) -- 2668
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(10,13)), 0, 10) -- 2669
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(12,15)), 0, 10) -- 2670
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(14,17)), 0, 10) -- 2671
,( 1, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(24,25),(16,19)), 0, 10) -- 2672
,( 1, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(26,27),(18,21)), 0, 10) -- 2673
,( 1, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(28,29),(20,23)), 0, 10) -- 2674
,( 1, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(30,31),(22,23)), 0, 10) -- 2675
,( 1, E,0,0,((24,25),(21,21),( 1, 1),(20,20),(23,23),(14,17)), 0, 10) -- 2676
,( 1, E,0,0,((26,27),(23,23),( 3, 3),(22,22),(25,25),(16,19)), 0, 10) -- 2677
,( 1, E,0,0,((28,29),(25,25),( 5, 5),(24,24),(27,27),(18,21)), 0, 10) -- 2678
,( 1, E,0,0,((30,31),(27,27),( 7, 7),(26,26),(29,29),(20,23)), 0, 10) -- 2679
,( 1, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(22,23),(16,19)), 0, 10) -- 2680
,( 1, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(24,25),(18,21)), 0, 10) -- 2681
,( 1, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(26,27),(20,23)), 0, 10) -- 2682
,( 1, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(28,29),(22,23)), 0, 10) -- 2683
,( 1, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 2684
,( 1, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 2685
,( 1, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 2686
,( 1, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 2687
,( 1, E,0,0,((22,25),(20,21),( 1, 1),(19,19),(24,24),(16,19)), 0, 10) -- 2688
,( 1, E,0,0,((24,27),(22,23),( 3, 3),(21,21),(26,26),(18,21)), 0, 10) -- 2689
,( 1, E,0,0,((26,29),(24,25),( 5, 5),(23,23),(28,28),(20,23)), 0, 10) -- 2690
,( 1, E,0,0,((28,31),(26,27),( 7, 7),(25,25),(30,30),(22,23)), 0, 10) -- 2691
,( 1, E,0,0,((24,25),(20,21),( 0, 1),(18,18),(19,19),( 6, 9)), 0, 10) -- 2692
,( 1, E,0,0,((26,27),(22,23),( 2, 3),(20,20),(21,21),( 8,11)), 0, 10) -- 2693
,( 1, E,0,0,((28,29),(24,25),( 4, 5),(22,22),(23,23),(10,13)), 0, 10) -- 2694
,( 1, E,0,0,((30,31),(26,27),( 6, 7),(24,24),(25,25),(12,15)), 0, 10) -- 2695
,( 1, E,0,0,((22,23),(20,20),( 0, 0),(18,18),(21,21),(12,15)), 0, 10) -- 2696
,( 1, E,0,0,((24,25),(22,22),( 2, 2),(20,20),(23,23),(14,17)), 0, 10) -- 2697
,( 1, E,0,0,((26,27),(24,24),( 4, 4),(22,22),(25,25),(16,19)), 0, 10) -- 2698
,( 1, E,0,0,((28,29),(26,26),( 6, 6),(24,24),(27,27),(18,21)), 0, 10) -- 2699
,( 1, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 8,11)), 0,  9) -- 2700
,( 1, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(10,13)), 0,  9) -- 2701
,( 1, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(12,15)), 0,  9) -- 2702
,( 1, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(14,17)), 0,  9) -- 2703
,( 1, E,0,0,((18,21),(18,19),( 0, 1),(20,21),(24,25),(12,15)), 0,  9) -- 2704
,( 1, E,0,0,((20,23),(20,21),( 2, 3),(22,23),(26,27),(14,17)), 0,  9) -- 2705
,( 1, E,0,0,((22,25),(22,23),( 4, 5),(24,25),(28,29),(16,19)), 0,  9) -- 2706
,( 1, E,0,0,((24,27),(24,25),( 6, 7),(26,27),(30,31),(18,21)), 0,  9) -- 2707
,( 1, E,0,0,((20,23),(20,21),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 2708
,( 1, E,0,0,((22,25),(22,23),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 2709
,( 1, E,0,0,((24,27),(24,25),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 2710
,( 1, E,0,0,((26,29),(26,27),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 2711
,( 1, E,0,0,((18,21),(18,19),( 0, 1),(20,21),(22,23),( 6, 9)), 0,  9) -- 2712
,( 1, E,0,0,((20,23),(20,21),( 2, 3),(22,23),(24,25),( 8,11)), 0,  9) -- 2713
,( 1, E,0,0,((22,25),(22,23),( 4, 5),(24,25),(26,27),(10,13)), 0,  9) -- 2714
,( 1, E,0,0,((24,27),(24,25),( 6, 7),(26,27),(28,29),(12,15)), 0,  9) -- 2715
,( 1, E,0,0,((18,21),(18,19),( 0, 0),(18,19),(18,19),( 2, 5)), 0,  9) -- 2716
,( 1, E,0,0,((20,23),(20,21),( 2, 2),(20,21),(20,21),( 4, 7)), 0,  9) -- 2717
,( 1, E,0,0,((22,25),(22,23),( 4, 4),(22,23),(22,23),( 6, 9)), 0,  9) -- 2718
,( 1, E,0,0,((24,27),(24,25),( 6, 6),(24,25),(24,25),( 8,11)), 0,  9) -- 2719
,( 1, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),( 4, 7)), 0,  9) -- 2720
,( 1, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),( 6, 9)), 0,  9) -- 2721
,( 1, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),( 8,11)), 0,  9) -- 2722
,( 1, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),(10,13)), 0,  9) -- 2723
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 2724
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 2725
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 2726
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 2727
,( 1, E,0,0,((18,21),(18,19),( 0, 1),(19,19),(22,23),( 6, 7)), 0,  9) -- 2728
,( 1, E,0,0,((20,23),(20,21),( 2, 3),(21,21),(24,25),( 8, 9)), 0,  9) -- 2729
,( 1, E,0,0,((22,25),(22,23),( 4, 5),(23,23),(26,27),(10,11)), 0,  9) -- 2730
,( 1, E,0,0,((24,27),(24,25),( 6, 7),(25,25),(28,29),(12,13)), 0,  9) -- 2731
,( 1, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(12,15)), 0,  9) -- 2732
,( 1, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(14,17)), 0,  9) -- 2733
,( 1, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(16,19)), 0,  9) -- 2734
,( 1, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(18,21)), 0,  9) -- 2735
,( 1, E,0,0,((20,23),(18,19),( 0, 1),(19,19),(24,24),(12,15)), 0,  9) -- 2736
,( 1, E,0,0,((22,25),(20,21),( 2, 3),(21,21),(26,26),(14,17)), 0,  9) -- 2737
,( 1, E,0,0,((24,27),(22,23),( 4, 5),(23,23),(28,28),(16,19)), 0,  9) -- 2738
,( 1, E,0,0,((26,29),(24,25),( 6, 7),(25,25),(30,30),(18,21)), 0,  9) -- 2739
,( 1, E,0,0,((20,23),(19,19),( 0, 0),(17,17),(18,19),( 2, 5)), 0,  9) -- 2740
,( 1, E,0,0,((22,25),(21,21),( 2, 2),(19,19),(20,21),( 4, 7)), 0,  9) -- 2741
,( 1, E,0,0,((24,27),(23,23),( 4, 4),(21,21),(22,23),( 6, 9)), 0,  9) -- 2742
,( 1, E,0,0,((26,29),(25,25),( 6, 6),(23,23),(24,25),( 8,11)), 0,  9) -- 2743
,( 1, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(20,21),(10,13)), 0,  9) -- 2744
,( 1, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(22,23),(12,15)), 0,  9) -- 2745
,( 1, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(24,25),(14,17)), 0,  9) -- 2746
,( 1, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(26,27),(16,19)), 0,  9) -- 2747
,( 1, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 2748
,( 1, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 2749
,( 1, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 2750
,( 1, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 2751
,( 1, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(24,25),(12,15)), 0,  9) -- 2752
,( 1, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(26,27),(14,17)), 0,  9) -- 2753
,( 1, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(28,29),(16,19)), 0,  9) -- 2754
,( 1, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(30,31),(18,21)), 0,  9) -- 2755
,( 1, E,0,0,((16,19),(17,17),( 0, 0),(18,19),(20,21),( 4, 7)), 0,  9) -- 2756
,( 1, E,0,0,((18,21),(19,19),( 2, 2),(20,21),(22,23),( 6, 9)), 0,  9) -- 2757
,( 1, E,0,0,((20,23),(21,21),( 4, 4),(22,23),(24,25),( 8,11)), 0,  9) -- 2758
,( 1, E,0,0,((22,25),(23,23),( 6, 6),(24,25),(26,27),(10,13)), 0,  9) -- 2759
,( 1, E,0,0,((18,19),(17,17),( 0, 0),(19,19),(22,23),( 6, 9)), 0,  9) -- 2760
,( 1, E,0,0,((20,21),(19,19),( 2, 2),(21,21),(24,25),( 8,11)), 0,  9) -- 2761
,( 1, E,0,0,((22,23),(21,21),( 4, 4),(23,23),(26,27),(10,13)), 0,  9) -- 2762
,( 1, E,0,0,((24,25),(23,23),( 6, 6),(25,25),(28,29),(12,15)), 0,  9) -- 2763
,( 1, E,0,0,((20,21),(18,18),( 0, 0),(18,19),(21,21),(10,13)), 0,  9) -- 2764
,( 1, E,0,0,((22,23),(20,20),( 2, 2),(20,21),(23,23),(12,15)), 0,  9) -- 2765
,( 1, E,0,0,((24,25),(22,22),( 4, 4),(22,23),(25,25),(14,17)), 0,  9) -- 2766
,( 1, E,0,0,((26,27),(24,24),( 6, 6),(24,25),(27,27),(16,19)), 0,  9) -- 2767
,( 1, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 2768
,( 1, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 2769
,( 1, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 2770
,( 1, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 2771
,( 1, E,0,0,((22,23),(19,19),( 0, 0),(17,17),(20,20),( 8,11)), 0,  9) -- 2772
,( 1, E,0,0,((24,25),(21,21),( 2, 2),(19,19),(22,22),(10,13)), 0,  9) -- 2773
,( 1, E,0,0,((26,27),(23,23),( 4, 4),(21,21),(24,24),(12,15)), 0,  9) -- 2774
,( 1, E,0,0,((28,29),(25,25),( 6, 6),(23,23),(26,26),(14,17)), 0,  9) -- 2775
,( 1, E,0,0,((20,23),(18,19),( 0, 1),(20,21),(24,25),(14,17)), 0,  9) -- 2776
,( 1, E,0,0,((22,25),(20,21),( 2, 3),(22,23),(26,27),(16,19)), 0,  9) -- 2777
,( 1, E,0,0,((24,27),(22,23),( 4, 5),(24,25),(28,29),(18,21)), 0,  9) -- 2778
,( 1, E,0,0,((26,29),(24,25),( 6, 7),(26,27),(30,31),(20,23)), 0,  9) -- 2779
,( 1, E,0,0,((20,23),(20,20),( 0, 1),(18,19),(18,19),( 6, 9)), 0,  9) -- 2780
,( 1, E,0,0,((22,25),(22,22),( 2, 3),(20,21),(20,21),( 8,11)), 0,  9) -- 2781
,( 1, E,0,0,((24,27),(24,24),( 4, 5),(22,23),(22,23),(10,13)), 0,  9) -- 2782
,( 1, E,0,0,((26,29),(26,26),( 6, 7),(24,25),(24,25),(12,15)), 0,  9) -- 2783
,( 1, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(22,25),(10,13)), 0,  8) -- 2784
,( 1, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(24,27),(12,15)), 0,  8) -- 2785
,( 1, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(26,29),(14,17)), 0,  8) -- 2786
,( 1, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(28,31),(16,19)), 0,  8) -- 2787
,( 1, E,0,0,((18,21),(18,21),( 0, 1),(18,21),(18,21),( 2, 5)), 0,  8) -- 2788
,( 1, E,0,0,((20,23),(20,23),( 2, 3),(20,23),(20,23),( 4, 7)), 0,  8) -- 2789
,( 1, E,0,0,((22,25),(22,25),( 4, 5),(22,25),(22,25),( 6, 9)), 0,  8) -- 2790
,( 1, E,0,0,((24,27),(24,27),( 6, 7),(24,27),(24,27),( 8,11)), 0,  8) -- 2791
,( 1, E,0,0,((18,21),(18,21),( 0, 1),(16,19),(16,19),(99,99)), 0,  8) -- 2792
,( 1, E,0,0,((20,23),(20,23),( 2, 3),(18,21),(18,21),(99,99)), 0,  8) -- 2793
,( 1, E,0,0,((22,25),(22,25),( 4, 5),(20,23),(20,23),(99,99)), 0,  8) -- 2794
,( 1, E,0,0,((24,27),(24,27),( 6, 7),(22,25),(22,25),(99,99)), 0,  8) -- 2795
,( 1, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(18,21),(99,99)), 0,  7) -- 2796
,( 1, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(20,23),(99,99)), 0,  7) -- 2797
,( 1, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(22,25),(99,99)), 0,  7) -- 2798
,( 1, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(24,27),(99,99)), 0,  7) -- 2799
,( 1, E,0,0,((16,19),(16,19),( 0, 1),(16,19),(14,17),(99,99)), 0,  7) -- 2800
,( 1, E,0,0,((18,21),(18,21),( 2, 3),(18,21),(16,19),(99,99)), 0,  7) -- 2801
,( 1, E,0,0,((20,23),(20,23),( 4, 5),(20,23),(18,21),(99,99)), 0,  7) -- 2802
,( 1, E,0,0,((22,25),(22,25),( 6, 7),(22,25),(20,23),(99,99)), 0,  7) -- 2803
,( 1, E,0,0,((12,15),(14,17),( 0, 1),(20,21),(22,25),(99,99)), 0,  7) -- 2804
,( 1, E,0,0,((14,17),(16,19),( 2, 3),(22,23),(24,27),(99,99)), 0,  7) -- 2805
,( 1, E,0,0,((16,19),(18,21),( 4, 5),(24,25),(26,29),(99,99)), 0,  7) -- 2806
,( 1, E,0,0,((18,21),(20,23),( 6, 7),(26,27),(28,31),(99,99)), 0,  7) -- 2807
,( 1, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 2808
,( 1, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 2809
,( 1, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 2810
,( 1, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 2811
,( 1, E,0,1,((14,17),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  7) -- 2812
,( 1, E,0,1,((16,19),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  7) -- 2813
,( 1, E,0,1,((18,21),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  7) -- 2814
,( 1, E,0,1,((20,23),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  7) -- 2815
,( 1, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 2816
,( 1, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 2817
,( 1, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 2818
,( 1, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 2819
,( 1, E,0,1,(( 8,11),(12,15),( 0, 1),(18,21),(99,99),(99,99)), 0,  6) -- 2820
,( 1, E,0,1,((10,13),(14,17),( 2, 3),(20,23),(99,99),(99,99)), 0,  6) -- 2821
,( 1, E,0,1,((12,15),(16,19),( 4, 5),(22,25),(99,99),(99,99)), 0,  6) -- 2822
,( 1, E,0,1,((14,17),(18,21),( 6, 7),(24,27),(99,99),(99,99)), 0,  6) -- 2823
,( 1, E,0,1,((10,13),(14,17),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 2824
,( 1, E,0,1,((12,15),(16,19),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 2825
,( 1, E,0,1,((14,17),(18,21),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 2826
,( 1, E,0,1,((16,19),(20,23),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 2827
,( 1, E,0,1,((16,17),(99,99),( 0, 1),(12,13),(99,99),(99,99)), 0,  5) -- 2828
,( 1, E,0,1,((18,19),(99,99),( 2, 3),(14,15),(99,99),(99,99)), 0,  5) -- 2829
,( 1, E,0,1,((20,21),(99,99),( 4, 5),(16,17),(99,99),(99,99)), 0,  5) -- 2830
,( 1, E,0,1,((22,23),(99,99),( 6, 7),(18,19),(99,99),(99,99)), 0,  5) -- 2831
,( 1, E,0,1,((20,23),(22,23),( 0, 1),(99,99),(99,99),(99,99)), 0,  5) -- 2832
,( 1, E,0,1,((22,25),(24,25),( 2, 3),(99,99),(99,99),(99,99)), 0,  5) -- 2833
,( 1, E,0,1,((24,27),(26,27),( 4, 5),(99,99),(99,99),(99,99)), 0,  5) -- 2834
,( 1, E,0,1,((26,29),(28,29),( 6, 7),(99,99),(99,99),(99,99)), 0,  5) -- 2835
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 2836
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 2837
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 2838
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 2839
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 2840
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 2841
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 2842
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 2843
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 2844
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 2845
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 2846
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 2847
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 2848
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 2849
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 2850
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 2851
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 2852
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 2853
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 2854
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 2855
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 2856
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 2857
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 2858
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 2859
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 2860
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 2861
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 2862
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 2863
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 2864
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 2865
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 2866
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 2867
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 30) -- 2868
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 30) -- 2869
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 30) -- 2870
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 30) -- 2871
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 30) -- 2872
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 30) -- 2873
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 30) -- 2874
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 30) -- 2875
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 30) -- 2876
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 30) -- 2877
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 30) -- 2878
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 30) -- 2879
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 30) -- 2880
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 30) -- 2881
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 30) -- 2882
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 30) -- 2883
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 30) -- 2884
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 30) -- 2885
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 30) -- 2886
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 30) -- 2887
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 30) -- 2888
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 30) -- 2889
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 30) -- 2890
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 30) -- 2891
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 29) -- 2892
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 29) -- 2893
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 29) -- 2894
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 29) -- 2895
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 29) -- 2896
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 29) -- 2897
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 29) -- 2898
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 29) -- 2899
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 29) -- 2900
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 29) -- 2901
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 29) -- 2902
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 29) -- 2903
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 29) -- 2904
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 29) -- 2905
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 29) -- 2906
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 29) -- 2907
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 28) -- 2908
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 28) -- 2909
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 28) -- 2910
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 28) -- 2911
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 28) -- 2912
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 28) -- 2913
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 28) -- 2914
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 28) -- 2915
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 27) -- 2916
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 27) -- 2917
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 27) -- 2918
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 27) -- 2919
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 27) -- 2920
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 27) -- 2921
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 27) -- 2922
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 27) -- 2923
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 25) -- 2924
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 25) -- 2925
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 25) -- 2926
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 25) -- 2927
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 25) -- 2928
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 25) -- 2929
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 25) -- 2930
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 25) -- 2931
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 25) -- 2932
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 25) -- 2933
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 25) -- 2934
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 25) -- 2935
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 25) -- 2936
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 25) -- 2937
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 25) -- 2938
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 25) -- 2939
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 24) -- 2940
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 24) -- 2941
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 24) -- 2942
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 24) -- 2943
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 24) -- 2944
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 24) -- 2945
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 24) -- 2946
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 24) -- 2947
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 23) -- 2948
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 23) -- 2949
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 23) -- 2950
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 23) -- 2951
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 23) -- 2952
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 23) -- 2953
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 23) -- 2954
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 23) -- 2955
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 21) -- 2956
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 21) -- 2957
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 21) -- 2958
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(19,19),(18,18),(10,10)), 1, 21) -- 2959
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(20,20),(19,19),(11,11)), 1, 21) -- 2960
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(21,21),(20,20),(12,12)), 1, 21) -- 2961
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(22,22),(21,21),(13,13)), 1, 21) -- 2962
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(23,23),(22,22),(14,14)), 1, 21) -- 2963
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 21) -- 2964
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 21) -- 2965
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 21) -- 2966
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 21) -- 2967
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 21) -- 2968
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 21) -- 2969
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 21) -- 2970
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 21) -- 2971
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 20) -- 2972
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 20) -- 2973
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 20) -- 2974
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 20) -- 2975
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 20) -- 2976
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 20) -- 2977
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 20) -- 2978
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 20) -- 2979
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 20) -- 2980
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 20) -- 2981
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 20) -- 2982
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 20) -- 2983
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 20) -- 2984
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 20) -- 2985
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 20) -- 2986
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 20) -- 2987
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 20) -- 2988
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 20) -- 2989
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 20) -- 2990
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(19,19),(19,19),(10,10)), 1, 20) -- 2991
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(20,20),(20,20),(11,11)), 1, 20) -- 2992
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(21,21),(21,21),(12,12)), 1, 20) -- 2993
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(22,22),(22,22),(13,13)), 1, 20) -- 2994
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(23,23),(23,23),(14,14)), 1, 20) -- 2995
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 20) -- 2996
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 20) -- 2997
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 20) -- 2998
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 20) -- 2999
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 20) -- 3000
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 20) -- 3001
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 20) -- 3002
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 20) -- 3003
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 3004
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 3005
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 3006
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 3007
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 3008
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 3009
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 3010
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 3011
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 3012
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 3013
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 3014
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 3015
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 3016
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 3017
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 3018
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 3019
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 3020
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 3021
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 3022
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 3023
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 3024
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 3025
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 3026
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 3027
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 3028
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 3029
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 3030
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 3031
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 3032
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 3033
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 3034
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 3035
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 3036
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 3037
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 3038
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 3039
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 3040
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 3041
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 3042
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 3043
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 3044
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 3045
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 3046
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 3047
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 3048
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 3049
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 3050
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 3051
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 3052
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 3053
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 3054
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 3055
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 3056
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 3057
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 3058
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 3059
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 3060
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 3061
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 3062
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 3063
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 3064
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 3065
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 3066
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 3067
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 18) -- 3068
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 18) -- 3069
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 18) -- 3070
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 18) -- 3071
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 18) -- 3072
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 18) -- 3073
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 18) -- 3074
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 18) -- 3075
,( 2, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 3076
,( 2, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 3077
,( 2, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 3078
,( 2, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 3079
,( 2, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 3080
,( 2, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 3081
,( 2, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 3082
,( 2, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 3083
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 3084
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 3085
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 3086
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 3087
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 3088
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 3089
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 3090
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 3091
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 3092
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 3093
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 3094
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 3095
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 3096
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 3097
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 3098
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 3099
,( 2, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 3100
,( 2, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 3101
,( 2, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 3102
,( 2, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 3103
,( 2, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 3104
,( 2, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 3105
,( 2, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 3106
,( 2, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 3107
,( 2, E,0,0,((34,34),(26,26),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 16) -- 3108
,( 2, E,0,0,((35,35),(27,27),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 16) -- 3109
,( 2, E,0,0,((36,36),(28,28),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 16) -- 3110
,( 2, E,0,0,((37,37),(29,29),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 16) -- 3111
,( 2, E,0,0,((38,38),(30,30),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 16) -- 3112
,( 2, E,0,0,((39,39),(31,31),( 5, 5),(19,19),(19,19),(10,10)), 1, 16) -- 3113
,( 2, E,0,0,((40,40),(32,32),( 6, 6),(20,20),(20,20),(11,11)), 1, 16) -- 3114
,( 2, E,0,0,((41,41),(33,33),( 7, 7),(21,21),(21,21),(12,12)), 1, 16) -- 3115
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 16) -- 3116
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 16) -- 3117
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 16) -- 3118
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 16) -- 3119
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 16) -- 3120
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 16) -- 3121
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 16) -- 3122
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 16) -- 3123
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 16) -- 3124
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 16) -- 3125
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 16) -- 3126
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 16) -- 3127
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 16) -- 3128
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 16) -- 3129
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 16) -- 3130
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 16) -- 3131
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 16) -- 3132
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 16) -- 3133
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 16) -- 3134
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 16) -- 3135
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 16) -- 3136
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 16) -- 3137
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 16) -- 3138
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 16) -- 3139
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 3140
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 3141
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 3142
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 3143
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 3144
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 3145
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 3146
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 3147
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 15) -- 3148
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 15) -- 3149
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 15) -- 3150
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 15) -- 3151
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 15) -- 3152
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),(10,10)), 1, 15) -- 3153
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(11,11)), 1, 15) -- 3154
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(12,12)), 1, 15) -- 3155
,( 2, E,0,0,((36,36),(27,27),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 3156
,( 2, E,0,0,((37,37),(28,28),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 3157
,( 2, E,0,0,((38,38),(29,29),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 3158
,( 2, E,0,0,((39,39),(30,30),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 3159
,( 2, E,0,0,((40,40),(31,31),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 3160
,( 2, E,0,0,((41,41),(32,32),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 3161
,( 2, E,0,0,((42,42),(33,33),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 3162
,( 2, E,0,0,((43,43),(34,34),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 3163
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 3, 3)), 1, 15) -- 3164
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 4, 4)), 1, 15) -- 3165
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 5, 5)), 1, 15) -- 3166
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 6, 6)), 1, 15) -- 3167
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 7, 7)), 1, 15) -- 3168
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 8, 8)), 1, 15) -- 3169
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),( 9, 9)), 1, 15) -- 3170
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(10,10)), 1, 15) -- 3171
,( 2, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 3172
,( 2, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 3173
,( 2, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 3174
,( 2, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 3175
,( 2, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 3176
,( 2, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 3177
,( 2, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 3178
,( 2, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 3179
,( 2, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 3180
,( 2, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 3181
,( 2, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 3182
,( 2, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 3183
,( 2, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 3184
,( 2, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 3185
,( 2, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 3186
,( 2, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 3187
,( 2, E,0,0,((36,36),(27,27),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 3188
,( 2, E,0,0,((37,37),(28,28),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 3189
,( 2, E,0,0,((38,38),(29,29),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 3190
,( 2, E,0,0,((39,39),(30,30),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 3191
,( 2, E,0,0,((40,40),(31,31),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 3192
,( 2, E,0,0,((41,41),(32,32),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 3193
,( 2, E,0,0,((42,42),(33,33),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 3194
,( 2, E,0,0,((43,43),(34,34),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 3195
,( 2, E,0,0,((36,36),(27,27),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 3196
,( 2, E,0,0,((37,37),(28,28),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 3197
,( 2, E,0,0,((38,38),(29,29),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 3198
,( 2, E,0,0,((39,39),(30,30),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 3199
,( 2, E,0,0,((40,40),(31,31),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 3200
,( 2, E,0,0,((41,41),(32,32),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 3201
,( 2, E,0,0,((42,42),(33,33),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 3202
,( 2, E,0,0,((43,43),(34,34),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 3203
,( 2, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 3204
,( 2, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 3205
,( 2, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 3206
,( 2, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 3207
,( 2, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 3208
,( 2, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 3209
,( 2, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 3210
,( 2, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 3211
,( 2, E,0,0,((36,39),(28,29),( 0, 1),(15,15),(14,15),( 4, 7)), 1, 14) -- 3212
,( 2, E,0,0,((38,41),(30,31),( 2, 3),(17,17),(16,17),( 6, 9)), 1, 14) -- 3213
,( 2, E,0,0,((40,43),(32,33),( 4, 5),(19,19),(18,19),( 8,11)), 1, 14) -- 3214
,( 2, E,0,0,((42,45),(34,35),( 6, 7),(21,21),(20,21),(10,13)), 1, 14) -- 3215
,( 2, E,0,0,((36,39),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 13) -- 3216
,( 2, E,0,0,((38,41),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 13) -- 3217
,( 2, E,0,0,((40,43),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 13) -- 3218
,( 2, E,0,0,((42,45),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 13) -- 3219
,( 2, E,0,0,((36,39),(28,29),( 1, 1),(16,16),(14,15),( 6, 9)), 1, 13) -- 3220
,( 2, E,0,0,((38,41),(30,31),( 3, 3),(18,18),(16,17),( 8,11)), 1, 13) -- 3221
,( 2, E,0,0,((40,43),(32,33),( 5, 5),(20,20),(18,19),(10,13)), 1, 13) -- 3222
,( 2, E,0,0,((42,45),(34,35),( 7, 7),(22,22),(20,21),(12,15)), 1, 13) -- 3223
,( 2, E,0,0,((36,39),(26,27),( 0, 0),(14,14),(12,13),( 4, 7)), 1, 12) -- 3224
,( 2, E,0,0,((38,41),(28,29),( 2, 2),(16,16),(14,15),( 6, 9)), 1, 12) -- 3225
,( 2, E,0,0,((40,43),(30,31),( 4, 4),(18,18),(16,17),( 8,11)), 1, 12) -- 3226
,( 2, E,0,0,((42,45),(32,33),( 6, 6),(20,20),(18,19),(10,13)), 1, 12) -- 3227
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(13,13),( 4, 7)), 1, 12) -- 3228
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(15,15),( 6, 9)), 1, 12) -- 3229
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(17,17),( 8,11)), 1, 12) -- 3230
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(19,19),(10,13)), 1, 12) -- 3231
,( 2, E,0,0,((36,39),(27,27),( 0, 0),(14,14),(12,13),( 0, 3)), 1, 12) -- 3232
,( 2, E,0,0,((38,41),(29,29),( 2, 2),(16,16),(14,15),( 2, 5)), 1, 12) -- 3233
,( 2, E,0,0,((40,43),(31,31),( 4, 4),(18,18),(16,17),( 4, 7)), 1, 12) -- 3234
,( 2, E,0,0,((42,45),(33,33),( 6, 6),(20,20),(18,19),( 6, 9)), 1, 12) -- 3235
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 12) -- 3236
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 8,11)), 1, 12) -- 3237
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(10,13)), 1, 12) -- 3238
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(12,15)), 1, 12) -- 3239
,( 2, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,12),( 0, 3)), 1, 12) -- 3240
,( 2, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,14),( 2, 5)), 1, 12) -- 3241
,( 2, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,16),( 4, 7)), 1, 12) -- 3242
,( 2, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,18),( 6, 9)), 1, 12) -- 3243
,( 2, E,0,0,((38,41),(28,29),( 0, 0),(12,13),(10,11),( 0, 3)), 1, 11) -- 3244
,( 2, E,0,0,((40,43),(30,31),( 2, 2),(14,15),(12,13),( 2, 5)), 1, 11) -- 3245
,( 2, E,0,0,((42,45),(32,33),( 4, 4),(16,17),(14,15),( 4, 7)), 1, 11) -- 3246
,( 2, E,0,0,((44,47),(34,35),( 6, 6),(18,19),(16,17),( 6, 9)), 1, 11) -- 3247
,( 2, E,0,0,((40,41),(29,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 3248
,( 2, E,0,0,((42,43),(31,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 3249
,( 2, E,0,0,((44,45),(33,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 3250
,( 2, E,0,0,((46,47),(35,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 3251
,( 2, E,0,0,((40,43),(30,31),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 3252
,( 2, E,0,0,((42,45),(32,33),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 3253
,( 2, E,0,0,((44,47),(34,35),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 3254
,( 2, E,0,0,((46,49),(36,37),( 6, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 3255
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(10,11),( 0, 3)), 1, 11) -- 3256
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(12,13),( 2, 5)), 1, 11) -- 3257
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(14,15),( 4, 7)), 1, 11) -- 3258
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(16,17),( 6, 9)), 1, 11) -- 3259
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 3260
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 3261
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 3262
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 3263
,( 2, E,0,0,((38,39),(28,28),( 0, 0),(13,13),(12,12),( 4, 7)), 1, 11) -- 3264
,( 2, E,0,0,((40,41),(30,30),( 2, 2),(15,15),(14,14),( 6, 9)), 1, 11) -- 3265
,( 2, E,0,0,((42,43),(32,32),( 4, 4),(17,17),(16,16),( 8,11)), 1, 11) -- 3266
,( 2, E,0,0,((44,45),(34,34),( 6, 6),(19,19),(18,18),(10,13)), 1, 11) -- 3267
,( 2, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,13),( 4, 7)), 1, 11) -- 3268
,( 2, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,15),( 6, 9)), 1, 11) -- 3269
,( 2, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,17),( 8,11)), 1, 11) -- 3270
,( 2, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,19),(10,13)), 1, 11) -- 3271
,( 2, E,0,0,((38,38),(27,27),( 0, 0),(13,13),(11,11),( 2, 5)), 1, 11) -- 3272
,( 2, E,0,0,((40,40),(29,29),( 2, 2),(15,15),(13,13),( 4, 7)), 1, 11) -- 3273
,( 2, E,0,0,((42,42),(31,31),( 4, 4),(17,17),(15,15),( 6, 9)), 1, 11) -- 3274
,( 2, E,0,0,((44,44),(33,33),( 6, 6),(19,19),(17,17),( 8,11)), 1, 11) -- 3275
,( 2, E,0,0,((40,41),(30,30),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 11) -- 3276
,( 2, E,0,0,((42,43),(32,32),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 11) -- 3277
,( 2, E,0,0,((44,45),(34,34),( 5, 5),(20,20),(18,19),( 8,11)), 1, 11) -- 3278
,( 2, E,0,0,((46,47),(36,36),( 7, 7),(22,22),(20,21),(10,13)), 1, 11) -- 3279
,( 2, E,0,0,((40,43),(30,31),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 3280
,( 2, E,0,0,((42,45),(32,33),( 2, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 3281
,( 2, E,0,0,((44,47),(34,35),( 4, 5),(18,19),(16,17),(10,13)), 1, 10) -- 3282
,( 2, E,0,0,((46,49),(36,37),( 6, 7),(20,21),(18,19),(12,15)), 1, 10) -- 3283
,( 2, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(10,11),( 4, 7)), 1, 10) -- 3284
,( 2, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(12,13),( 6, 9)), 1, 10) -- 3285
,( 2, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(14,15),( 8,11)), 1, 10) -- 3286
,( 2, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(16,17),(10,13)), 1, 10) -- 3287
,( 2, E,0,0,((40,43),(30,31),( 0, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 3288
,( 2, E,0,0,((42,45),(32,33),( 2, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 3289
,( 2, E,0,0,((44,47),(34,35),( 4, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 3290
,( 2, E,0,0,((46,49),(36,37),( 6, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 3291
,( 2, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),( 6, 9)), 1, 10) -- 3292
,( 2, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),( 8,11)), 1, 10) -- 3293
,( 2, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),(10,13)), 1, 10) -- 3294
,( 2, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),(12,15)), 1, 10) -- 3295
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1, 10) -- 3296
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1, 10) -- 3297
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1, 10) -- 3298
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1, 10) -- 3299
,( 2, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(14,14),( 6, 9)), 1, 10) -- 3300
,( 2, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(16,16),( 8,11)), 1, 10) -- 3301
,( 2, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(18,18),(10,13)), 1, 10) -- 3302
,( 2, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(20,20),(12,15)), 1, 10) -- 3303
,( 2, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 10) -- 3304
,( 2, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 10) -- 3305
,( 2, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 10) -- 3306
,( 2, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,18),( 8,11)), 1, 10) -- 3307
,( 2, E,0,0,((40,43),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 1)), 1, 10) -- 3308
,( 2, E,0,0,((42,45),(32,33),( 2, 3),(14,15),(10,11),( 2, 3)), 1, 10) -- 3309
,( 2, E,0,0,((44,47),(34,35),( 4, 5),(16,17),(12,13),( 4, 5)), 1, 10) -- 3310
,( 2, E,0,0,((46,49),(36,37),( 6, 7),(18,19),(14,15),( 6, 7)), 1, 10) -- 3311
,( 2, E,0,0,((40,43),(30,31),( 0, 1),(14,14),(10,11),( 0, 1)), 1, 10) -- 3312
,( 2, E,0,0,((42,45),(32,33),( 2, 3),(16,16),(12,13),( 2, 3)), 1, 10) -- 3313
,( 2, E,0,0,((44,47),(34,35),( 4, 5),(18,18),(14,15),( 4, 5)), 1, 10) -- 3314
,( 2, E,0,0,((46,49),(36,37),( 6, 7),(20,20),(16,17),( 6, 7)), 1, 10) -- 3315
,( 2, E,0,0,((40,43),(30,30),( 0, 1),(12,13),(10,11),( 2, 5)), 1, 10) -- 3316
,( 2, E,0,0,((42,45),(32,32),( 2, 3),(14,15),(12,13),( 4, 7)), 1, 10) -- 3317
,( 2, E,0,0,((44,47),(34,34),( 4, 5),(16,17),(14,15),( 6, 9)), 1, 10) -- 3318
,( 2, E,0,0,((46,49),(36,36),( 6, 7),(18,19),(16,17),( 8,11)), 1, 10) -- 3319
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 3320
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 3321
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(10,13)), 1,  9) -- 3322
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(12,15)), 1,  9) -- 3323
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),(10,13)), 1,  9) -- 3324
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(12,15)), 1,  9) -- 3325
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(14,17)), 1,  9) -- 3326
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(16,19)), 1,  9) -- 3327
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 6, 9)), 1,  9) -- 3328
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),( 8,11)), 1,  9) -- 3329
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(10,13)), 1,  9) -- 3330
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(12,15)), 1,  9) -- 3331
,( 2, E,0,0,((40,43),(29,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1,  9) -- 3332
,( 2, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(12,13),( 8,11)), 1,  9) -- 3333
,( 2, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(14,15),(10,13)), 1,  9) -- 3334
,( 2, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(16,17),(12,15)), 1,  9) -- 3335
,( 2, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 4, 7)), 1,  9) -- 3336
,( 2, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 6, 9)), 1,  9) -- 3337
,( 2, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 8,11)), 1,  9) -- 3338
,( 2, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),(10,13)), 1,  9) -- 3339
,( 2, E,0,0,((40,43),(30,31),( 1, 1),(14,15),(14,15),(12,15)), 1,  9) -- 3340
,( 2, E,0,0,((42,45),(32,33),( 3, 3),(16,17),(16,17),(14,17)), 1,  9) -- 3341
,( 2, E,0,0,((44,47),(34,35),( 5, 5),(18,19),(18,19),(16,19)), 1,  9) -- 3342
,( 2, E,0,0,((46,49),(36,37),( 7, 7),(20,21),(20,21),(18,21)), 1,  9) -- 3343
,( 2, E,0,0,((40,43),(29,29),( 0, 1),(14,15),(14,15),(14,17)), 1,  9) -- 3344
,( 2, E,0,0,((42,45),(31,31),( 2, 3),(16,17),(16,17),(16,19)), 1,  9) -- 3345
,( 2, E,0,0,((44,47),(33,33),( 4, 5),(18,19),(18,19),(18,21)), 1,  9) -- 3346
,( 2, E,0,0,((46,49),(35,35),( 6, 7),(20,21),(20,21),(20,23)), 1,  9) -- 3347
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 2, 5)), 1,  9) -- 3348
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 4, 7)), 1,  9) -- 3349
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 6, 9)), 1,  9) -- 3350
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 8,11)), 1,  9) -- 3351
,( 2, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),(10,13)), 1,  9) -- 3352
,( 2, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),(12,15)), 1,  9) -- 3353
,( 2, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(14,17)), 1,  9) -- 3354
,( 2, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(16,19)), 1,  9) -- 3355
,( 2, E,0,0,((42,45),(31,31),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 3356
,( 2, E,0,0,((44,47),(33,33),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 3357
,( 2, E,0,0,((46,49),(35,35),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 3358
,( 2, E,0,0,((48,51),(37,37),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 3359
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),(10,13)), 1,  9) -- 3360
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),(12,15)), 1,  9) -- 3361
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(14,17)), 1,  9) -- 3362
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(16,19)), 1,  9) -- 3363
,( 2, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(12,13),(10,13)), 1,  9) -- 3364
,( 2, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(14,15),(12,15)), 1,  9) -- 3365
,( 2, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(16,17),(14,17)), 1,  9) -- 3366
,( 2, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(18,19),(16,19)), 1,  9) -- 3367
,( 2, E,0,0,((40,43),(29,29),( 0, 0),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 3368
,( 2, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(10,11),( 2, 5)), 1,  9) -- 3369
,( 2, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(12,13),( 4, 7)), 1,  9) -- 3370
,( 2, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(14,15),( 6, 9)), 1,  9) -- 3371
,( 2, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(11,11),(10,13)), 1,  9) -- 3372
,( 2, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(13,13),(12,15)), 1,  9) -- 3373
,( 2, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(15,15),(14,17)), 1,  9) -- 3374
,( 2, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(17,17),(16,19)), 1,  9) -- 3375
,( 2, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),(14,17)), 1,  9) -- 3376
,( 2, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(16,19)), 1,  9) -- 3377
,( 2, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(18,21)), 1,  9) -- 3378
,( 2, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(20,23)), 1,  9) -- 3379
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,14),(13,13),(14,17)), 1,  9) -- 3380
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,16),(15,15),(16,19)), 1,  9) -- 3381
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,18),(17,17),(18,21)), 1,  9) -- 3382
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,20),(19,19),(20,23)), 1,  9) -- 3383
,( 2, E,0,0,((44,47),(32,33),( 1, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 3384
,( 2, E,0,0,((46,49),(34,35),( 3, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 3385
,( 2, E,0,0,((48,51),(36,37),( 5, 5),(16,17),(14,15),(10,13)), 1,  9) -- 3386
,( 2, E,0,0,((50,53),(38,39),( 7, 7),(18,19),(16,17),(12,15)), 1,  9) -- 3387
,( 2, E,0,0,((44,47),(32,32),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 3388
,( 2, E,0,0,((46,49),(34,34),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 3389
,( 2, E,0,0,((48,51),(36,36),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 3390
,( 2, E,0,0,((50,53),(38,38),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 3391
,( 2, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(14,15),(17,17)), 1,  9) -- 3392
,( 2, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(16,17),(19,19)), 1,  9) -- 3393
,( 2, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(18,19),(21,21)), 1,  9) -- 3394
,( 2, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(20,21),(23,23)), 1,  9) -- 3395
,( 2, E,0,0,((44,45),(32,32),( 1, 1),(14,14),(12,13),( 6, 9)), 1,  9) -- 3396
,( 2, E,0,0,((46,47),(34,34),( 3, 3),(16,16),(14,15),( 8,11)), 1,  9) -- 3397
,( 2, E,0,0,((48,49),(36,36),( 5, 5),(18,18),(16,17),(10,13)), 1,  9) -- 3398
,( 2, E,0,0,((50,51),(38,38),( 7, 7),(20,20),(18,19),(12,15)), 1,  9) -- 3399
,( 2, E,0,0,((40,43),(29,29),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 3400
,( 2, E,0,0,((42,45),(31,31),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 3401
,( 2, E,0,0,((44,47),(33,33),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 3402
,( 2, E,0,0,((46,49),(35,35),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 3403
,( 2, E,0,0,((42,45),(32,32),( 1, 1),(14,14),(10,11),( 4, 7)), 1,  9) -- 3404
,( 2, E,0,0,((44,47),(34,34),( 3, 3),(16,16),(12,13),( 6, 9)), 1,  9) -- 3405
,( 2, E,0,0,((46,49),(36,36),( 5, 5),(18,18),(14,15),( 8,11)), 1,  9) -- 3406
,( 2, E,0,0,((48,51),(38,38),( 7, 7),(20,20),(16,17),(10,13)), 1,  9) -- 3407
,( 2, E,0,0,((44,44),(31,31),( 1, 1),(14,14),(12,13),( 6, 9)), 1,  9) -- 3408
,( 2, E,0,0,((46,46),(33,33),( 3, 3),(16,16),(14,15),( 8,11)), 1,  9) -- 3409
,( 2, E,0,0,((48,48),(35,35),( 5, 5),(18,18),(16,17),(10,13)), 1,  9) -- 3410
,( 2, E,0,0,((50,50),(37,37),( 7, 7),(20,20),(18,19),(12,15)), 1,  9) -- 3411
,( 2, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(16,16),(14,14)), 1,  9) -- 3412
,( 2, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(18,18),(16,16)), 1,  9) -- 3413
,( 2, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(20,20),(18,18)), 1,  9) -- 3414
,( 2, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(22,22),(20,20)), 1,  9) -- 3415
,( 2, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),(12,15)), 1,  9) -- 3416
,( 2, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),(14,17)), 1,  9) -- 3417
,( 2, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),(16,19)), 1,  9) -- 3418
,( 2, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),(18,21)), 1,  9) -- 3419
,( 2, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(12,15),(11,11)), 1,  8) -- 3420
,( 2, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(14,17),(13,13)), 1,  8) -- 3421
,( 2, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(16,19),(15,15)), 1,  8) -- 3422
,( 2, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(18,21),(17,17)), 1,  8) -- 3423
,( 2, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 8,11),( 6, 9)), 1,  8) -- 3424
,( 2, E,0,0,((46,49),(32,35),( 2, 3),(12,15),(10,13),( 8,11)), 1,  8) -- 3425
,( 2, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(12,15),(10,13)), 1,  8) -- 3426
,( 2, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(14,17),(12,15)), 1,  8) -- 3427
,( 2, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 3428
,( 2, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 3429
,( 2, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 3430
,( 2, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 3431
,( 2, E,0,0,((46,49),(32,35),( 0, 1),(12,15),(10,13),(99,99)), 1,  7) -- 3432
,( 2, E,0,0,((48,51),(34,37),( 2, 3),(14,17),(12,15),(99,99)), 1,  7) -- 3433
,( 2, E,0,0,((50,53),(36,39),( 4, 5),(16,19),(14,17),(99,99)), 1,  7) -- 3434
,( 2, E,0,0,((52,55),(38,41),( 6, 7),(18,21),(16,19),(99,99)), 1,  7) -- 3435
,( 2, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(16,19),(99,99)), 1,  7) -- 3436
,( 2, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(18,21),(99,99)), 1,  7) -- 3437
,( 2, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(20,23),(99,99)), 1,  7) -- 3438
,( 2, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(22,25),(99,99)), 1,  7) -- 3439
,( 2, E,0,1,((48,51),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 3440
,( 2, E,0,1,((50,53),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 3441
,( 2, E,0,1,((52,55),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 3442
,( 2, E,0,1,((54,57),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 3443
,( 2, E,0,1,((44,47),(30,33),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 3444
,( 2, E,0,1,((46,49),(32,35),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 3445
,( 2, E,0,1,((48,51),(34,37),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 3446
,( 2, E,0,1,((50,53),(36,39),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 3447
,( 2, E,0,1,((42,45),(28,31),( 0, 1),(16,17),(99,99),(99,99)), 1,  6) -- 3448
,( 2, E,0,1,((44,47),(30,33),( 2, 3),(18,19),(99,99),(99,99)), 1,  6) -- 3449
,( 2, E,0,1,((46,49),(32,35),( 4, 5),(20,21),(99,99),(99,99)), 1,  6) -- 3450
,( 2, E,0,1,((48,51),(34,37),( 6, 7),(22,23),(99,99),(99,99)), 1,  6) -- 3451
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 3452
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 3453
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 3454
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 3455
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 3456
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 3457
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 3458
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 3459
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 3460
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 3461
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 3462
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 3463
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 3464
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 3465
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 3466
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 3467
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 3468
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 3469
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 3470
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 3471
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 3472
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 3473
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 3474
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 3475
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 3476
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 3477
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 3478
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 3479
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 3480
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 3481
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 3482
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 3483
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 3484
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 3485
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 3486
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 3487
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 3488
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 3489
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 3490
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 3491
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 3492
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 3493
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 3494
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 3495
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 3496
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 3497
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 3498
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 3499
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 3500
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 3501
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 3502
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 3503
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 3504
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 3505
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 3506
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 3507
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 30) -- 3508
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 30) -- 3509
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 30) -- 3510
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 30) -- 3511
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 30) -- 3512
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 30) -- 3513
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 30) -- 3514
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 30) -- 3515
,( 2, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 30) -- 3516
,( 2, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 30) -- 3517
,( 2, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 0, 30) -- 3518
,( 2, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 0, 30) -- 3519
,( 2, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 0, 30) -- 3520
,( 2, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 0, 30) -- 3521
,( 2, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 0, 30) -- 3522
,( 2, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 0, 30) -- 3523
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 29) -- 3524
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 29) -- 3525
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 29) -- 3526
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 29) -- 3527
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 29) -- 3528
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 29) -- 3529
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 29) -- 3530
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 29) -- 3531
,( 2, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 29) -- 3532
,( 2, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 29) -- 3533
,( 2, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 29) -- 3534
,( 2, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 29) -- 3535
,( 2, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 29) -- 3536
,( 2, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 29) -- 3537
,( 2, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 29) -- 3538
,( 2, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 29) -- 3539
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 26) -- 3540
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 26) -- 3541
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 26) -- 3542
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 26) -- 3543
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 26) -- 3544
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 26) -- 3545
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 26) -- 3546
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 26) -- 3547
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 24) -- 3548
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 24) -- 3549
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 24) -- 3550
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 24) -- 3551
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 24) -- 3552
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 24) -- 3553
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 24) -- 3554
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 24) -- 3555
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 23) -- 3556
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 23) -- 3557
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 23) -- 3558
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 23) -- 3559
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 23) -- 3560
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 23) -- 3561
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 23) -- 3562
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 23) -- 3563
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 23) -- 3564
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 23) -- 3565
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 23) -- 3566
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 23) -- 3567
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 23) -- 3568
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 23) -- 3569
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 23) -- 3570
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 23) -- 3571
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 22) -- 3572
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 22) -- 3573
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 22) -- 3574
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 22) -- 3575
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 22) -- 3576
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 22) -- 3577
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 22) -- 3578
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 22) -- 3579
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 22) -- 3580
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 22) -- 3581
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 22) -- 3582
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 22) -- 3583
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 22) -- 3584
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 22) -- 3585
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 22) -- 3586
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 22) -- 3587
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 21) -- 3588
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 21) -- 3589
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 21) -- 3590
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 21) -- 3591
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 21) -- 3592
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 21) -- 3593
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 21) -- 3594
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 21) -- 3595
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 21) -- 3596
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 21) -- 3597
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 21) -- 3598
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 21) -- 3599
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 21) -- 3600
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 21) -- 3601
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 21) -- 3602
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 21) -- 3603
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 20) -- 3604
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 20) -- 3605
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 20) -- 3606
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 20) -- 3607
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 20) -- 3608
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 20) -- 3609
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 20) -- 3610
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 20) -- 3611
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 3612
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 3613
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 3614
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 3615
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 3616
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 3617
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 3618
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 3619
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 19) -- 3620
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 19) -- 3621
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 19) -- 3622
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 19) -- 3623
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 19) -- 3624
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 19) -- 3625
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 19) -- 3626
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 19) -- 3627
,( 2, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 3628
,( 2, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 3629
,( 2, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 3630
,( 2, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 3631
,( 2, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 3632
,( 2, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 3633
,( 2, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 3634
,( 2, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 3635
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 3636
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 3637
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 3638
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 3639
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 3640
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 3641
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 3642
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 3643
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 3644
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 3645
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 3646
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 3647
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 3648
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 3649
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 3650
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 3651
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 3652
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 3653
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 3654
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 3655
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 3656
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 3657
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 3658
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 3659
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 18) -- 3660
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 18) -- 3661
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 18) -- 3662
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 18) -- 3663
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 18) -- 3664
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 18) -- 3665
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 18) -- 3666
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 18) -- 3667
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 18) -- 3668
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 18) -- 3669
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 18) -- 3670
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 18) -- 3671
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 18) -- 3672
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 18) -- 3673
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 18) -- 3674
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 18) -- 3675
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 18) -- 3676
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 18) -- 3677
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 18) -- 3678
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 18) -- 3679
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 18) -- 3680
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 18) -- 3681
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 18) -- 3682
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 18) -- 3683
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 17) -- 3684
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 17) -- 3685
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 17) -- 3686
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 17) -- 3687
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 17) -- 3688
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 17) -- 3689
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 17) -- 3690
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 17) -- 3691
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 3692
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 3693
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 3694
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 3695
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 3696
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 3697
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 3698
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 3699
,( 2, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 3700
,( 2, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 3701
,( 2, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 3702
,( 2, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 3703
,( 2, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 3704
,( 2, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 3705
,( 2, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 3706
,( 2, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 3707
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 16) -- 3708
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 16) -- 3709
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 16) -- 3710
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 16) -- 3711
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 16) -- 3712
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 16) -- 3713
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 16) -- 3714
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 16) -- 3715
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 16) -- 3716
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 16) -- 3717
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 16) -- 3718
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 16) -- 3719
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 16) -- 3720
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 16) -- 3721
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 16) -- 3722
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 16) -- 3723
,( 2, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 3724
,( 2, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 3725
,( 2, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 3726
,( 2, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 3727
,( 2, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 3728
,( 2, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 3729
,( 2, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 3730
,( 2, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 3731
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(12,12)), 0, 16) -- 3732
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(13,13)), 0, 16) -- 3733
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(14,14)), 0, 16) -- 3734
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(15,15)), 0, 16) -- 3735
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(16,16)), 0, 16) -- 3736
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(17,17)), 0, 16) -- 3737
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(18,18)), 0, 16) -- 3738
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(19,19)), 0, 16) -- 3739
,( 2, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 16) -- 3740
,( 2, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 16) -- 3741
,( 2, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 16) -- 3742
,( 2, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 16) -- 3743
,( 2, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 16) -- 3744
,( 2, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 16) -- 3745
,( 2, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 16) -- 3746
,( 2, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 16) -- 3747
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 3748
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 3749
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 3750
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 3751
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 3752
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 3753
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 3754
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 3755
,( 2, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),( 9, 9)), 0, 16) -- 3756
,( 2, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(10,10)), 0, 16) -- 3757
,( 2, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(11,11)), 0, 16) -- 3758
,( 2, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(12,12)), 0, 16) -- 3759
,( 2, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(13,13)), 0, 16) -- 3760
,( 2, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(14,14)), 0, 16) -- 3761
,( 2, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(15,15)), 0, 16) -- 3762
,( 2, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(16,16)), 0, 16) -- 3763
,( 2, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 15) -- 3764
,( 2, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 15) -- 3765
,( 2, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 15) -- 3766
,( 2, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 15) -- 3767
,( 2, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 15) -- 3768
,( 2, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 15) -- 3769
,( 2, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 15) -- 3770
,( 2, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 15) -- 3771
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 3772
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 3773
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 3774
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 3775
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 3776
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 3777
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 3778
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 3779
,( 2, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 15) -- 3780
,( 2, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 15) -- 3781
,( 2, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 15) -- 3782
,( 2, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 15) -- 3783
,( 2, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 15) -- 3784
,( 2, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 15) -- 3785
,( 2, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 15) -- 3786
,( 2, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 15) -- 3787
,( 2, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 15) -- 3788
,( 2, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 15) -- 3789
,( 2, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 15) -- 3790
,( 2, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 15) -- 3791
,( 2, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 15) -- 3792
,( 2, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 15) -- 3793
,( 2, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 15) -- 3794
,( 2, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 15) -- 3795
,( 2, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 15) -- 3796
,( 2, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 15) -- 3797
,( 2, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 15) -- 3798
,( 2, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 15) -- 3799
,( 2, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 15) -- 3800
,( 2, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 15) -- 3801
,( 2, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 15) -- 3802
,( 2, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 15) -- 3803
,( 2, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 3804
,( 2, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 3805
,( 2, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 3806
,( 2, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 3807
,( 2, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 3808
,( 2, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 3809
,( 2, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 3810
,( 2, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 3811
,( 2, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 3812
,( 2, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 3813
,( 2, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 3814
,( 2, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 3815
,( 2, E,0,0,((28,31),(24,24),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 3816
,( 2, E,0,0,((30,33),(26,26),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 3817
,( 2, E,0,0,((32,35),(28,28),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 3818
,( 2, E,0,0,((34,37),(30,30),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 3819
,( 2, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(12,15)), 0, 14) -- 3820
,( 2, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(14,17)), 0, 14) -- 3821
,( 2, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(16,19)), 0, 14) -- 3822
,( 2, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(18,21)), 0, 14) -- 3823
,( 2, E,0,0,((26,27),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 13) -- 3824
,( 2, E,0,0,((28,29),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 13) -- 3825
,( 2, E,0,0,((30,31),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 13) -- 3826
,( 2, E,0,0,((32,33),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 13) -- 3827
,( 2, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),( 6, 9)), 0, 13) -- 3828
,( 2, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),( 8,11)), 0, 13) -- 3829
,( 2, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(10,13)), 0, 13) -- 3830
,( 2, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(12,15)), 0, 13) -- 3831
,( 2, E,0,0,((24,27),(20,21),( 0, 1),(17,17),(20,21),(12,15)), 0, 12) -- 3832
,( 2, E,0,0,((26,29),(22,23),( 2, 3),(19,19),(22,23),(14,17)), 0, 12) -- 3833
,( 2, E,0,0,((28,31),(24,25),( 4, 5),(21,21),(24,25),(16,19)), 0, 12) -- 3834
,( 2, E,0,0,((30,33),(26,27),( 6, 7),(23,23),(26,27),(18,21)), 0, 12) -- 3835
,( 2, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),( 8,11)), 0, 12) -- 3836
,( 2, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(10,13)), 0, 12) -- 3837
,( 2, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(12,15)), 0, 12) -- 3838
,( 2, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(14,17)), 0, 12) -- 3839
,( 2, E,0,0,((24,27),(21,21),( 0, 0),(17,17),(18,19),( 8,11)), 0, 12) -- 3840
,( 2, E,0,0,((26,29),(23,23),( 2, 2),(19,19),(20,21),(10,13)), 0, 12) -- 3841
,( 2, E,0,0,((28,31),(25,25),( 4, 4),(21,21),(22,23),(12,15)), 0, 12) -- 3842
,( 2, E,0,0,((30,33),(27,27),( 6, 6),(23,23),(24,25),(14,17)), 0, 12) -- 3843
,( 2, E,0,0,((26,29),(22,23),( 1, 1),(19,19),(22,23),(14,17)), 0, 12) -- 3844
,( 2, E,0,0,((28,31),(24,25),( 3, 3),(21,21),(24,25),(16,19)), 0, 12) -- 3845
,( 2, E,0,0,((30,33),(26,27),( 5, 5),(23,23),(26,27),(18,21)), 0, 12) -- 3846
,( 2, E,0,0,((32,35),(28,29),( 7, 7),(25,25),(28,29),(20,23)), 0, 12) -- 3847
,( 2, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(10,13)), 0, 12) -- 3848
,( 2, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(12,15)), 0, 12) -- 3849
,( 2, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(14,17)), 0, 12) -- 3850
,( 2, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(16,19)), 0, 12) -- 3851
,( 2, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(18,19),( 8,11)), 0, 12) -- 3852
,( 2, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(20,21),(10,13)), 0, 12) -- 3853
,( 2, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(22,23),(12,15)), 0, 12) -- 3854
,( 2, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(24,25),(14,17)), 0, 12) -- 3855
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 3856
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 3857
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 3858
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 3859
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(17,17),(18,19),( 8,11)), 0, 11) -- 3860
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(19,19),(20,21),(10,13)), 0, 11) -- 3861
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(21,21),(22,23),(12,15)), 0, 11) -- 3862
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(23,23),(24,25),(14,17)), 0, 11) -- 3863
,( 2, E,0,0,((24,27),(22,23),( 0, 1),(19,19),(22,23),(12,15)), 0, 11) -- 3864
,( 2, E,0,0,((26,29),(24,25),( 2, 3),(21,21),(24,25),(14,17)), 0, 11) -- 3865
,( 2, E,0,0,((28,31),(26,27),( 4, 5),(23,23),(26,27),(16,19)), 0, 11) -- 3866
,( 2, E,0,0,((30,33),(28,29),( 6, 7),(25,25),(28,29),(18,21)), 0, 11) -- 3867
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 11) -- 3868
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 11) -- 3869
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 11) -- 3870
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 11) -- 3871
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(10,13)), 0, 11) -- 3872
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(12,15)), 0, 11) -- 3873
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(14,17)), 0, 11) -- 3874
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(16,19)), 0, 11) -- 3875
,( 2, E,0,0,((24,27),(20,21),( 0, 1),(17,17),(18,19),( 4, 7)), 0, 11) -- 3876
,( 2, E,0,0,((26,29),(22,23),( 2, 3),(19,19),(20,21),( 6, 9)), 0, 11) -- 3877
,( 2, E,0,0,((28,31),(24,25),( 4, 5),(21,21),(22,23),( 8,11)), 0, 11) -- 3878
,( 2, E,0,0,((30,33),(26,27),( 6, 7),(23,23),(24,25),(10,13)), 0, 11) -- 3879
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(17,17),(20,21),( 8,11)), 0, 11) -- 3880
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(19,19),(22,23),(10,13)), 0, 11) -- 3881
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(21,21),(24,25),(12,15)), 0, 11) -- 3882
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(23,23),(26,27),(14,17)), 0, 11) -- 3883
,( 2, E,0,0,((25,25),(22,22),( 0, 1),(18,19),(20,21),(10,13)), 0, 11) -- 3884
,( 2, E,0,0,((27,27),(24,24),( 2, 3),(20,21),(22,23),(12,15)), 0, 11) -- 3885
,( 2, E,0,0,((29,29),(26,26),( 4, 5),(22,23),(24,25),(14,17)), 0, 11) -- 3886
,( 2, E,0,0,((31,31),(28,28),( 6, 7),(24,25),(26,27),(16,19)), 0, 11) -- 3887
,( 2, E,0,0,((26,29),(24,24),( 1, 1),(99,99),(22,23),(12,15)), 0, 11) -- 3888
,( 2, E,0,0,((28,31),(26,26),( 3, 3),(99,99),(24,25),(14,17)), 0, 11) -- 3889
,( 2, E,0,0,((30,33),(28,28),( 5, 5),(99,99),(26,27),(16,19)), 0, 11) -- 3890
,( 2, E,0,0,((32,35),(30,30),( 7, 7),(99,99),(28,29),(18,21)), 0, 11) -- 3891
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 3892
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 3893
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 3894
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 3895
,( 2, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),(10,13)), 0, 10) -- 3896
,( 2, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),(12,15)), 0, 10) -- 3897
,( 2, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(14,17)), 0, 10) -- 3898
,( 2, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(16,19)), 0, 10) -- 3899
,( 2, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 3900
,( 2, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 3901
,( 2, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 3902
,( 2, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 3903
,( 2, E,0,0,((22,23),(20,21),( 0, 1),(17,17),(18,19),( 4, 7)), 0, 10) -- 3904
,( 2, E,0,0,((24,25),(22,23),( 2, 3),(19,19),(20,21),( 6, 9)), 0, 10) -- 3905
,( 2, E,0,0,((26,27),(24,25),( 4, 5),(21,21),(22,23),( 8,11)), 0, 10) -- 3906
,( 2, E,0,0,((28,29),(26,27),( 6, 7),(23,23),(24,25),(10,13)), 0, 10) -- 3907
,( 2, E,0,0,((20,23),(18,19),( 0, 1),(17,17),(18,19),( 6, 9)), 0, 10) -- 3908
,( 2, E,0,0,((22,25),(20,21),( 2, 3),(19,19),(20,21),( 8,11)), 0, 10) -- 3909
,( 2, E,0,0,((24,27),(22,23),( 4, 5),(21,21),(22,23),(10,13)), 0, 10) -- 3910
,( 2, E,0,0,((26,29),(24,25),( 6, 7),(23,23),(24,25),(12,15)), 0, 10) -- 3911
,( 2, E,0,0,((20,23),(18,19),( 0, 0),(18,18),(20,21),( 6, 9)), 0, 10) -- 3912
,( 2, E,0,0,((22,25),(20,21),( 2, 2),(20,20),(22,23),( 8,11)), 0, 10) -- 3913
,( 2, E,0,0,((24,27),(22,23),( 4, 4),(22,22),(24,25),(10,13)), 0, 10) -- 3914
,( 2, E,0,0,((26,29),(24,25),( 6, 6),(24,24),(26,27),(12,15)), 0, 10) -- 3915
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 2, 5)), 0, 10) -- 3916
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 4, 7)), 0, 10) -- 3917
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),( 6, 9)), 0, 10) -- 3918
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),( 8,11)), 0, 10) -- 3919
,( 2, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 8,11)), 0, 10) -- 3920
,( 2, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(10,13)), 0, 10) -- 3921
,( 2, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(12,15)), 0, 10) -- 3922
,( 2, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(14,17)), 0, 10) -- 3923
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(19,19),(22,23),( 8, 9)), 0, 10) -- 3924
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(21,21),(24,25),(10,11)), 0, 10) -- 3925
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(23,23),(26,27),(12,13)), 0, 10) -- 3926
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(25,25),(28,29),(14,15)), 0, 10) -- 3927
,( 2, E,0,0,((24,27),(22,23),( 0, 1),(99,99),(20,21),( 6, 9)), 0, 10) -- 3928
,( 2, E,0,0,((26,29),(24,25),( 2, 3),(99,99),(22,23),( 8,11)), 0, 10) -- 3929
,( 2, E,0,0,((28,31),(26,27),( 4, 5),(99,99),(24,25),(10,13)), 0, 10) -- 3930
,( 2, E,0,0,((30,33),(28,29),( 6, 7),(99,99),(26,27),(12,15)), 0, 10) -- 3931
,( 2, E,0,0,((24,27),(22,22),( 0, 1),(99,99),(18,19),( 4, 7)), 0, 10) -- 3932
,( 2, E,0,0,((26,29),(24,24),( 2, 3),(99,99),(20,21),( 6, 9)), 0, 10) -- 3933
,( 2, E,0,0,((28,31),(26,26),( 4, 5),(99,99),(22,23),( 8,11)), 0, 10) -- 3934
,( 2, E,0,0,((30,33),(28,28),( 6, 7),(99,99),(24,25),(10,13)), 0, 10) -- 3935
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 3936
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 3937
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 3938
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 3939
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 0, 3)), 0,  9) -- 3940
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 2, 5)), 0,  9) -- 3941
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 4, 7)), 0,  9) -- 3942
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),( 6, 9)), 0,  9) -- 3943
,( 2, E,0,0,((20,23),(20,20),( 0, 1),(18,19),(20,21),( 8,11)), 0,  9) -- 3944
,( 2, E,0,0,((22,25),(22,22),( 2, 3),(20,21),(22,23),(10,13)), 0,  9) -- 3945
,( 2, E,0,0,((24,27),(24,24),( 4, 5),(22,23),(24,25),(12,15)), 0,  9) -- 3946
,( 2, E,0,0,((26,29),(26,26),( 6, 7),(24,25),(26,27),(14,17)), 0,  9) -- 3947
,( 2, E,0,0,((20,23),(20,21),( 1, 1),(20,20),(22,23),( 6, 9)), 0,  9) -- 3948
,( 2, E,0,0,((22,25),(22,23),( 3, 3),(22,22),(24,25),( 8,11)), 0,  9) -- 3949
,( 2, E,0,0,((24,27),(24,25),( 5, 5),(24,24),(26,27),(10,13)), 0,  9) -- 3950
,( 2, E,0,0,((26,29),(26,27),( 7, 7),(26,26),(28,29),(12,15)), 0,  9) -- 3951
,( 2, E,0,0,((20,23),(18,19),( 0, 1),(17,17),(18,19),( 0, 3)), 0,  9) -- 3952
,( 2, E,0,0,((22,25),(20,21),( 2, 3),(19,19),(20,21),( 2, 5)), 0,  9) -- 3953
,( 2, E,0,0,((24,27),(22,23),( 4, 5),(21,21),(22,23),( 4, 7)), 0,  9) -- 3954
,( 2, E,0,0,((26,29),(24,25),( 6, 7),(23,23),(24,25),( 6, 9)), 0,  9) -- 3955
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(20,20),(22,23),( 4, 7)), 0,  9) -- 3956
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(22,22),(24,25),( 6, 9)), 0,  9) -- 3957
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(24,24),(26,27),( 8,11)), 0,  9) -- 3958
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(26,26),(28,29),(10,13)), 0,  9) -- 3959
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(20,20),(24,25),(12,15)), 0,  9) -- 3960
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(22,22),(26,27),(14,17)), 0,  9) -- 3961
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(24,24),(28,29),(16,19)), 0,  9) -- 3962
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(26,26),(30,31),(18,21)), 0,  9) -- 3963
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 4, 7)), 0,  9) -- 3964
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 6, 9)), 0,  9) -- 3965
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 8,11)), 0,  9) -- 3966
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),(10,13)), 0,  9) -- 3967
,( 2, E,0,0,((16,19),(16,17),( 0, 1),(19,19),(22,23),( 3, 3)), 0,  9) -- 3968
,( 2, E,0,0,((18,21),(18,19),( 2, 3),(21,21),(24,25),( 5, 5)), 0,  9) -- 3969
,( 2, E,0,0,((20,23),(20,21),( 4, 5),(23,23),(26,27),( 7, 7)), 0,  9) -- 3970
,( 2, E,0,0,((22,25),(22,23),( 6, 7),(25,25),(28,29),( 9, 9)), 0,  9) -- 3971
,( 2, E,0,0,((20,23),(20,21),( 0, 1),(19,19),(22,23),( 2, 5)), 0,  9) -- 3972
,( 2, E,0,0,((22,25),(22,23),( 2, 3),(21,21),(24,25),( 4, 7)), 0,  9) -- 3973
,( 2, E,0,0,((24,27),(24,25),( 4, 5),(23,23),(26,27),( 6, 9)), 0,  9) -- 3974
,( 2, E,0,0,((26,29),(26,27),( 6, 7),(25,25),(28,29),( 8,11)), 0,  9) -- 3975
,( 2, E,0,0,((22,25),(20,21),( 1, 1),(19,19),(24,25),(14,17)), 0,  9) -- 3976
,( 2, E,0,0,((24,27),(22,23),( 3, 3),(21,21),(26,27),(16,19)), 0,  9) -- 3977
,( 2, E,0,0,((26,29),(24,25),( 5, 5),(23,23),(28,29),(18,21)), 0,  9) -- 3978
,( 2, E,0,0,((28,31),(26,27),( 7, 7),(25,25),(30,31),(20,23)), 0,  9) -- 3979
,( 2, E,0,0,((22,22),(19,19),( 0, 0),(18,18),(20,20),( 2, 5)), 0,  9) -- 3980
,( 2, E,0,0,((24,24),(21,21),( 2, 2),(20,20),(22,22),( 4, 7)), 0,  9) -- 3981
,( 2, E,0,0,((26,26),(23,23),( 4, 4),(22,22),(24,24),( 6, 9)), 0,  9) -- 3982
,( 2, E,0,0,((28,28),(25,25),( 6, 6),(24,24),(26,26),( 8,11)), 0,  9) -- 3983
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(18,18),(20,21),( 0, 1)), 0,  9) -- 3984
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(20,20),(22,23),( 2, 3)), 0,  9) -- 3985
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(22,22),(24,25),( 4, 5)), 0,  9) -- 3986
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(24,24),(26,27),( 6, 7)), 0,  9) -- 3987
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 3988
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 3989
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 3990
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 3991
,( 2, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(16,17),( 0, 1)), 0,  9) -- 3992
,( 2, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(18,19),( 2, 3)), 0,  9) -- 3993
,( 2, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(20,21),( 4, 5)), 0,  9) -- 3994
,( 2, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(22,23),( 6, 7)), 0,  9) -- 3995
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(17,17),(16,17),(99,99)), 0,  9) -- 3996
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(19,19),(18,19),(99,99)), 0,  9) -- 3997
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(21,21),(20,21),(99,99)), 0,  9) -- 3998
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(23,23),(22,23),(99,99)), 0,  9) -- 3999
,( 2, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(18,19),(99,99)), 0,  9) -- 4000
,( 2, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(20,21),(99,99)), 0,  9) -- 4001
,( 2, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(22,23),(99,99)), 0,  9) -- 4002
,( 2, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(24,25),(99,99)), 0,  9) -- 4003
,( 2, E,0,0,((24,25),(22,22),( 1, 1),(99,99),(20,21),( 2, 5)), 0,  9) -- 4004
,( 2, E,0,0,((26,27),(24,24),( 3, 3),(99,99),(22,23),( 4, 7)), 0,  9) -- 4005
,( 2, E,0,0,((28,29),(26,26),( 5, 5),(99,99),(24,25),( 6, 9)), 0,  9) -- 4006
,( 2, E,0,0,((30,31),(28,28),( 7, 7),(99,99),(26,27),( 8,11)), 0,  9) -- 4007
,( 2, E,0,0,((24,27),(22,23),( 1, 1),(99,99),(22,22),( 6, 9)), 0,  9) -- 4008
,( 2, E,0,0,((26,29),(24,25),( 3, 3),(99,99),(24,24),( 8,11)), 0,  9) -- 4009
,( 2, E,0,0,((28,31),(26,27),( 5, 5),(99,99),(26,26),(10,13)), 0,  9) -- 4010
,( 2, E,0,0,((30,33),(28,29),( 7, 7),(99,99),(28,28),(12,15)), 0,  9) -- 4011
,( 2, E,0,0,((16,19),(16,17),( 0, 0),(99,99),(21,21),(99,99)), 0,  9) -- 4012
,( 2, E,0,0,((18,21),(18,19),( 2, 2),(99,99),(23,23),(99,99)), 0,  9) -- 4013
,( 2, E,0,0,((20,23),(20,21),( 4, 4),(99,99),(25,25),(99,99)), 0,  9) -- 4014
,( 2, E,0,0,((22,25),(22,23),( 6, 6),(99,99),(27,27),(99,99)), 0,  9) -- 4015
,( 2, E,0,0,((16,19),(16,19),( 0, 1),(16,19),(18,21),(99,99)), 0,  8) -- 4016
,( 2, E,0,0,((18,21),(18,21),( 2, 3),(18,21),(20,23),(99,99)), 0,  8) -- 4017
,( 2, E,0,0,((20,23),(20,23),( 4, 5),(20,23),(22,25),(99,99)), 0,  8) -- 4018
,( 2, E,0,0,((22,25),(22,25),( 6, 7),(22,25),(24,27),(99,99)), 0,  8) -- 4019
,( 2, E,0,0,((18,21),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 4020
,( 2, E,0,0,((20,23),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 4021
,( 2, E,0,0,((22,25),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 4022
,( 2, E,0,0,((24,27),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 4023
,( 2, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(14,17),(99,99)), 0,  8) -- 4024
,( 2, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(16,19),(99,99)), 0,  8) -- 4025
,( 2, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(18,21),(99,99)), 0,  8) -- 4026
,( 2, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(20,23),(99,99)), 0,  8) -- 4027
,( 2, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(16,19),(99,99)), 0,  8) -- 4028
,( 2, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(18,21),(99,99)), 0,  8) -- 4029
,( 2, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(20,23),(99,99)), 0,  8) -- 4030
,( 2, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(22,25),(99,99)), 0,  8) -- 4031
,( 2, E,0,1,((16,19),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  7) -- 4032
,( 2, E,0,1,((18,21),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  7) -- 4033
,( 2, E,0,1,((20,23),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  7) -- 4034
,( 2, E,0,1,((22,25),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  7) -- 4035
,( 2, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 4036
,( 2, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 4037
,( 2, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 4038
,( 2, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 4039
,( 2, E,0,1,((20,23),(18,21),( 0, 1),(99,99),(99,99),(99,99)), 0,  7) -- 4040
,( 2, E,0,1,((22,25),(20,23),( 2, 3),(99,99),(99,99),(99,99)), 0,  7) -- 4041
,( 2, E,0,1,((24,27),(22,25),( 4, 5),(99,99),(99,99),(99,99)), 0,  7) -- 4042
,( 2, E,0,1,((26,29),(24,27),( 6, 7),(99,99),(99,99),(99,99)), 0,  7) -- 4043
,( 2, E,0,1,((12,15),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 4044
,( 2, E,0,1,((14,17),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 4045
,( 2, E,0,1,((16,19),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 4046
,( 2, E,0,1,((18,21),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 4047
,( 2, E,0,1,((18,21),(20,23),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 4048
,( 2, E,0,1,((20,23),(22,25),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 4049
,( 2, E,0,1,((22,25),(24,27),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 4050
,( 2, E,0,1,((24,27),(26,29),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 4051
,( 2, E,0,1,(( 8,11),(12,15),( 0, 1),(99,99),(99,99),(99,99)), 0,  6) -- 4052
,( 2, E,0,1,((10,13),(14,17),( 2, 3),(99,99),(99,99),(99,99)), 0,  6) -- 4053
,( 2, E,0,1,((12,15),(16,19),( 4, 5),(99,99),(99,99),(99,99)), 0,  6) -- 4054
,( 2, E,0,1,((14,17),(18,21),( 6, 7),(99,99),(99,99),(99,99)), 0,  6) -- 4055
,( 2, E,0,1,((16,17),(18,21),( 0, 1),(12,12),(99,99),(99,99)), 0,  5) -- 4056
,( 2, E,0,1,((18,19),(20,23),( 2, 3),(14,14),(99,99),(99,99)), 0,  5) -- 4057
,( 2, E,0,1,((20,21),(22,25),( 4, 5),(16,16),(99,99),(99,99)), 0,  5) -- 4058
,( 2, E,0,1,((22,23),(24,27),( 6, 7),(18,18),(99,99),(99,99)), 0,  5) -- 4059
,( 3, E,0,0,((32,32),(24,24),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 31) -- 4060
,( 3, E,0,0,((33,33),(25,25),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 31) -- 4061
,( 3, E,0,0,((34,34),(26,26),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 31) -- 4062
,( 3, E,0,0,((35,35),(27,27),( 3, 3),(99,99),(19,19),(10,10)), 1, 31) -- 4063
,( 3, E,0,0,((36,36),(28,28),( 4, 4),(99,99),(20,20),(11,11)), 1, 31) -- 4064
,( 3, E,0,0,((37,37),(29,29),( 5, 5),(99,99),(21,21),(12,12)), 1, 31) -- 4065
,( 3, E,0,0,((38,38),(30,30),( 6, 6),(99,99),(22,22),(13,13)), 1, 31) -- 4066
,( 3, E,0,0,((39,39),(31,31),( 7, 7),(99,99),(23,23),(14,14)), 1, 31) -- 4067
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(17,17),( 8, 8)), 1, 31) -- 4068
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(18,18),( 9, 9)), 1, 31) -- 4069
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(19,19),(10,10)), 1, 31) -- 4070
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(20,20),(11,11)), 1, 31) -- 4071
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(21,21),(12,12)), 1, 31) -- 4072
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(22,22),(13,13)), 1, 31) -- 4073
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(23,23),(14,14)), 1, 31) -- 4074
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(24,24),(15,15)), 1, 31) -- 4075
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(16,16),( 8, 8)), 1, 31) -- 4076
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(17,17),( 9, 9)), 1, 31) -- 4077
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(18,18),(10,10)), 1, 31) -- 4078
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(19,19),(11,11)), 1, 31) -- 4079
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(20,20),(12,12)), 1, 31) -- 4080
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(21,21),(13,13)), 1, 31) -- 4081
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(22,22),(14,14)), 1, 31) -- 4082
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(23,23),(15,15)), 1, 31) -- 4083
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 31) -- 4084
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 31) -- 4085
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 31) -- 4086
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(19,19),(10,10)), 1, 31) -- 4087
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(20,20),(11,11)), 1, 31) -- 4088
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(21,21),(12,12)), 1, 31) -- 4089
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(22,22),(13,13)), 1, 31) -- 4090
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(23,23),(14,14)), 1, 31) -- 4091
,( 3, E,0,0,((32,32),(24,24),( 0, 0),(99,99),(16,16),( 8, 8)), 1, 31) -- 4092
,( 3, E,0,0,((33,33),(25,25),( 1, 1),(99,99),(17,17),( 9, 9)), 1, 31) -- 4093
,( 3, E,0,0,((34,34),(26,26),( 2, 2),(99,99),(18,18),(10,10)), 1, 31) -- 4094
,( 3, E,0,0,((35,35),(27,27),( 3, 3),(99,99),(19,19),(11,11)), 1, 31) -- 4095
,( 3, E,0,0,((36,36),(28,28),( 4, 4),(99,99),(20,20),(12,12)), 1, 31) -- 4096
,( 3, E,0,0,((37,37),(29,29),( 5, 5),(99,99),(21,21),(13,13)), 1, 31) -- 4097
,( 3, E,0,0,((38,38),(30,30),( 6, 6),(99,99),(22,22),(14,14)), 1, 31) -- 4098
,( 3, E,0,0,((39,39),(31,31),( 7, 7),(99,99),(23,23),(15,15)), 1, 31) -- 4099
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 31) -- 4100
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 31) -- 4101
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 31) -- 4102
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(19,19),(10,10)), 1, 31) -- 4103
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(20,20),(11,11)), 1, 31) -- 4104
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(21,21),(12,12)), 1, 31) -- 4105
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(22,22),(13,13)), 1, 31) -- 4106
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(23,23),(14,14)), 1, 31) -- 4107
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(17,17),( 8, 8)), 1, 31) -- 4108
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(18,18),( 9, 9)), 1, 31) -- 4109
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(19,19),(10,10)), 1, 31) -- 4110
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(20,20),(11,11)), 1, 31) -- 4111
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(21,21),(12,12)), 1, 31) -- 4112
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(22,22),(13,13)), 1, 31) -- 4113
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(23,23),(14,14)), 1, 31) -- 4114
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(24,24),(15,15)), 1, 31) -- 4115
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 28) -- 4116
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 28) -- 4117
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 28) -- 4118
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(19,19),(10,10)), 1, 28) -- 4119
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(20,20),(11,11)), 1, 28) -- 4120
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(21,21),(12,12)), 1, 28) -- 4121
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(22,22),(13,13)), 1, 28) -- 4122
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(23,23),(14,14)), 1, 28) -- 4123
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(16,16),( 8, 8)), 1, 27) -- 4124
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(17,17),( 9, 9)), 1, 27) -- 4125
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(18,18),(10,10)), 1, 27) -- 4126
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(19,19),(11,11)), 1, 27) -- 4127
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(20,20),(12,12)), 1, 27) -- 4128
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(21,21),(13,13)), 1, 27) -- 4129
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(22,22),(14,14)), 1, 27) -- 4130
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(23,23),(15,15)), 1, 27) -- 4131
,( 3, E,0,0,((32,32),(24,24),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 24) -- 4132
,( 3, E,0,0,((33,33),(25,25),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 24) -- 4133
,( 3, E,0,0,((34,34),(26,26),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 24) -- 4134
,( 3, E,0,0,((35,35),(27,27),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 24) -- 4135
,( 3, E,0,0,((36,36),(28,28),( 4, 4),(99,99),(19,19),(10,10)), 1, 24) -- 4136
,( 3, E,0,0,((37,37),(29,29),( 5, 5),(99,99),(20,20),(11,11)), 1, 24) -- 4137
,( 3, E,0,0,((38,38),(30,30),( 6, 6),(99,99),(21,21),(12,12)), 1, 24) -- 4138
,( 3, E,0,0,((39,39),(31,31),( 7, 7),(99,99),(22,22),(13,13)), 1, 24) -- 4139
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 24) -- 4140
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 24) -- 4141
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 24) -- 4142
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 24) -- 4143
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(19,19),(10,10)), 1, 24) -- 4144
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(20,20),(11,11)), 1, 24) -- 4145
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(21,21),(12,12)), 1, 24) -- 4146
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(22,22),(13,13)), 1, 24) -- 4147
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(16,16),( 6, 6)), 1, 23) -- 4148
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(17,17),( 7, 7)), 1, 23) -- 4149
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(18,18),( 8, 8)), 1, 23) -- 4150
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(19,19),( 9, 9)), 1, 23) -- 4151
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(20,20),(10,10)), 1, 23) -- 4152
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(21,21),(11,11)), 1, 23) -- 4153
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(22,22),(12,12)), 1, 23) -- 4154
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(23,23),(13,13)), 1, 23) -- 4155
,( 3, E,0,0,((33,33),(26,26),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 23) -- 4156
,( 3, E,0,0,((34,34),(27,27),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 23) -- 4157
,( 3, E,0,0,((35,35),(28,28),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 23) -- 4158
,( 3, E,0,0,((36,36),(29,29),( 3, 3),(99,99),(19,19),(10,10)), 1, 23) -- 4159
,( 3, E,0,0,((37,37),(30,30),( 4, 4),(99,99),(20,20),(11,11)), 1, 23) -- 4160
,( 3, E,0,0,((38,38),(31,31),( 5, 5),(99,99),(21,21),(12,12)), 1, 23) -- 4161
,( 3, E,0,0,((39,39),(32,32),( 6, 6),(99,99),(22,22),(13,13)), 1, 23) -- 4162
,( 3, E,0,0,((40,40),(33,33),( 7, 7),(99,99),(23,23),(14,14)), 1, 23) -- 4163
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 23) -- 4164
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 23) -- 4165
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 23) -- 4166
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 23) -- 4167
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(19,19),(10,10)), 1, 23) -- 4168
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(20,20),(11,11)), 1, 23) -- 4169
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(21,21),(12,12)), 1, 23) -- 4170
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(22,22),(13,13)), 1, 23) -- 4171
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(15,15),( 7, 7)), 1, 22) -- 4172
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(16,16),( 8, 8)), 1, 22) -- 4173
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(17,17),( 9, 9)), 1, 22) -- 4174
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(18,18),(10,10)), 1, 22) -- 4175
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(19,19),(11,11)), 1, 22) -- 4176
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(20,20),(12,12)), 1, 22) -- 4177
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(21,21),(13,13)), 1, 22) -- 4178
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(22,22),(14,14)), 1, 22) -- 4179
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 21) -- 4180
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 21) -- 4181
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 21) -- 4182
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(19,19),(10,10)), 1, 21) -- 4183
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(20,20),(11,11)), 1, 21) -- 4184
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(21,21),(12,12)), 1, 21) -- 4185
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(22,22),(13,13)), 1, 21) -- 4186
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(23,23),(14,14)), 1, 21) -- 4187
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(16,16),( 6, 6)), 1, 20) -- 4188
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(17,17),( 7, 7)), 1, 20) -- 4189
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(18,18),( 8, 8)), 1, 20) -- 4190
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(19,19),( 9, 9)), 1, 20) -- 4191
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(20,20),(10,10)), 1, 20) -- 4192
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(21,21),(11,11)), 1, 20) -- 4193
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(22,22),(12,12)), 1, 20) -- 4194
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(23,23),(13,13)), 1, 20) -- 4195
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 19) -- 4196
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 19) -- 4197
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 19) -- 4198
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 19) -- 4199
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(19,19),(10,10)), 1, 19) -- 4200
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(20,20),(11,11)), 1, 19) -- 4201
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(21,21),(12,12)), 1, 19) -- 4202
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(22,22),(13,13)), 1, 19) -- 4203
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 19) -- 4204
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 19) -- 4205
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 19) -- 4206
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 19) -- 4207
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(19,19),(10,10)), 1, 19) -- 4208
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(20,20),(11,11)), 1, 19) -- 4209
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(21,21),(12,12)), 1, 19) -- 4210
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(22,22),(13,13)), 1, 19) -- 4211
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(16,16),( 7, 7)), 1, 19) -- 4212
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(17,17),( 8, 8)), 1, 19) -- 4213
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(18,18),( 9, 9)), 1, 19) -- 4214
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(19,19),(10,10)), 1, 19) -- 4215
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(20,20),(11,11)), 1, 19) -- 4216
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(21,21),(12,12)), 1, 19) -- 4217
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(22,22),(13,13)), 1, 19) -- 4218
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(23,23),(14,14)), 1, 19) -- 4219
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(15,15),( 6, 6)), 1, 18) -- 4220
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(16,16),( 7, 7)), 1, 18) -- 4221
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(17,17),( 8, 8)), 1, 18) -- 4222
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(18,18),( 9, 9)), 1, 18) -- 4223
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(19,19),(10,10)), 1, 18) -- 4224
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(20,20),(11,11)), 1, 18) -- 4225
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(21,21),(12,12)), 1, 18) -- 4226
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(22,22),(13,13)), 1, 18) -- 4227
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(15,15),( 5, 5)), 1, 18) -- 4228
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(16,16),( 6, 6)), 1, 18) -- 4229
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(17,17),( 7, 7)), 1, 18) -- 4230
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(18,18),( 8, 8)), 1, 18) -- 4231
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(19,19),( 9, 9)), 1, 18) -- 4232
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(20,20),(10,10)), 1, 18) -- 4233
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(21,21),(11,11)), 1, 18) -- 4234
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(22,22),(12,12)), 1, 18) -- 4235
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(15,15),( 5, 5)), 1, 18) -- 4236
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(16,16),( 6, 6)), 1, 18) -- 4237
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(17,17),( 7, 7)), 1, 18) -- 4238
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(18,18),( 8, 8)), 1, 18) -- 4239
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(19,19),( 9, 9)), 1, 18) -- 4240
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(20,20),(10,10)), 1, 18) -- 4241
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(21,21),(11,11)), 1, 18) -- 4242
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(22,22),(12,12)), 1, 18) -- 4243
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(15,15),( 7, 7)), 1, 18) -- 4244
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(16,16),( 8, 8)), 1, 18) -- 4245
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(17,17),( 9, 9)), 1, 18) -- 4246
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(18,18),(10,10)), 1, 18) -- 4247
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(19,19),(11,11)), 1, 18) -- 4248
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(20,20),(12,12)), 1, 18) -- 4249
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(21,21),(13,13)), 1, 18) -- 4250
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(22,22),(14,14)), 1, 18) -- 4251
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(15,15),( 7, 7)), 1, 18) -- 4252
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(16,16),( 8, 8)), 1, 18) -- 4253
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(17,17),( 9, 9)), 1, 18) -- 4254
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(18,18),(10,10)), 1, 18) -- 4255
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(19,19),(11,11)), 1, 18) -- 4256
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(20,20),(12,12)), 1, 18) -- 4257
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(21,21),(13,13)), 1, 18) -- 4258
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(22,22),(14,14)), 1, 18) -- 4259
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(15,15),( 5, 5)), 1, 17) -- 4260
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(16,16),( 6, 6)), 1, 17) -- 4261
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(17,17),( 7, 7)), 1, 17) -- 4262
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(18,18),( 8, 8)), 1, 17) -- 4263
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(19,19),( 9, 9)), 1, 17) -- 4264
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(20,20),(10,10)), 1, 17) -- 4265
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(21,21),(11,11)), 1, 17) -- 4266
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(22,22),(12,12)), 1, 17) -- 4267
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(14,14),( 5, 5)), 1, 17) -- 4268
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(15,15),( 6, 6)), 1, 17) -- 4269
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(16,16),( 7, 7)), 1, 17) -- 4270
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(17,17),( 8, 8)), 1, 17) -- 4271
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(18,18),( 9, 9)), 1, 17) -- 4272
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(19,19),(10,10)), 1, 17) -- 4273
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(20,20),(11,11)), 1, 17) -- 4274
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(21,21),(12,12)), 1, 17) -- 4275
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(14,14),( 6, 6)), 1, 17) -- 4276
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(15,15),( 7, 7)), 1, 17) -- 4277
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(16,16),( 8, 8)), 1, 17) -- 4278
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(17,17),( 9, 9)), 1, 17) -- 4279
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(18,18),(10,10)), 1, 17) -- 4280
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(19,19),(11,11)), 1, 17) -- 4281
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(20,20),(12,12)), 1, 17) -- 4282
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(21,21),(13,13)), 1, 17) -- 4283
,( 3, E,0,0,((33,33),(25,25),( 0, 0),(99,99),(14,14),( 5, 5)), 1, 17) -- 4284
,( 3, E,0,0,((34,34),(26,26),( 1, 1),(99,99),(15,15),( 6, 6)), 1, 17) -- 4285
,( 3, E,0,0,((35,35),(27,27),( 2, 2),(99,99),(16,16),( 7, 7)), 1, 17) -- 4286
,( 3, E,0,0,((36,36),(28,28),( 3, 3),(99,99),(17,17),( 8, 8)), 1, 17) -- 4287
,( 3, E,0,0,((37,37),(29,29),( 4, 4),(99,99),(18,18),( 9, 9)), 1, 17) -- 4288
,( 3, E,0,0,((38,38),(30,30),( 5, 5),(99,99),(19,19),(10,10)), 1, 17) -- 4289
,( 3, E,0,0,((39,39),(31,31),( 6, 6),(99,99),(20,20),(11,11)), 1, 17) -- 4290
,( 3, E,0,0,((40,40),(32,32),( 7, 7),(99,99),(21,21),(12,12)), 1, 17) -- 4291
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(14,14),( 6, 6)), 1, 17) -- 4292
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(15,15),( 7, 7)), 1, 17) -- 4293
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(16,16),( 8, 8)), 1, 17) -- 4294
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(17,17),( 9, 9)), 1, 17) -- 4295
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(18,18),(10,10)), 1, 17) -- 4296
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(19,19),(11,11)), 1, 17) -- 4297
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(20,20),(12,12)), 1, 17) -- 4298
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(21,21),(13,13)), 1, 17) -- 4299
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(14,14),( 5, 5)), 1, 17) -- 4300
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(15,15),( 6, 6)), 1, 17) -- 4301
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(16,16),( 7, 7)), 1, 17) -- 4302
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(17,17),( 8, 8)), 1, 17) -- 4303
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(18,18),( 9, 9)), 1, 17) -- 4304
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(19,19),(10,10)), 1, 17) -- 4305
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(20,20),(11,11)), 1, 17) -- 4306
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(21,21),(12,12)), 1, 17) -- 4307
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(14,14),( 5, 5)), 1, 16) -- 4308
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(15,15),( 6, 6)), 1, 16) -- 4309
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(16,16),( 7, 7)), 1, 16) -- 4310
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(17,17),( 8, 8)), 1, 16) -- 4311
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(18,18),( 9, 9)), 1, 16) -- 4312
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(19,19),(10,10)), 1, 16) -- 4313
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(20,20),(11,11)), 1, 16) -- 4314
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(21,21),(12,12)), 1, 16) -- 4315
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(14,14),( 4, 4)), 1, 16) -- 4316
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(15,15),( 5, 5)), 1, 16) -- 4317
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(16,16),( 6, 6)), 1, 16) -- 4318
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(17,17),( 7, 7)), 1, 16) -- 4319
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(18,18),( 8, 8)), 1, 16) -- 4320
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(19,19),( 9, 9)), 1, 16) -- 4321
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(20,20),(10,10)), 1, 16) -- 4322
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(21,21),(11,11)), 1, 16) -- 4323
,( 3, E,0,0,((34,34),(26,26),( 0, 0),(99,99),(14,14),( 4, 4)), 1, 16) -- 4324
,( 3, E,0,0,((35,35),(27,27),( 1, 1),(99,99),(15,15),( 5, 5)), 1, 16) -- 4325
,( 3, E,0,0,((36,36),(28,28),( 2, 2),(99,99),(16,16),( 6, 6)), 1, 16) -- 4326
,( 3, E,0,0,((37,37),(29,29),( 3, 3),(99,99),(17,17),( 7, 7)), 1, 16) -- 4327
,( 3, E,0,0,((38,38),(30,30),( 4, 4),(99,99),(18,18),( 8, 8)), 1, 16) -- 4328
,( 3, E,0,0,((39,39),(31,31),( 5, 5),(99,99),(19,19),( 9, 9)), 1, 16) -- 4329
,( 3, E,0,0,((40,40),(32,32),( 6, 6),(99,99),(20,20),(10,10)), 1, 16) -- 4330
,( 3, E,0,0,((41,41),(33,33),( 7, 7),(99,99),(21,21),(11,11)), 1, 16) -- 4331
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(13,13),( 4, 4)), 1, 15) -- 4332
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(14,14),( 5, 5)), 1, 15) -- 4333
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(15,15),( 6, 6)), 1, 15) -- 4334
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(16,16),( 7, 7)), 1, 15) -- 4335
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(17,17),( 8, 8)), 1, 15) -- 4336
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(18,18),( 9, 9)), 1, 15) -- 4337
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(19,19),(10,10)), 1, 15) -- 4338
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(20,20),(11,11)), 1, 15) -- 4339
,( 3, E,0,0,((36,36),(27,27),( 0, 0),(99,99),(14,14),( 4, 4)), 1, 15) -- 4340
,( 3, E,0,0,((37,37),(28,28),( 1, 1),(99,99),(15,15),( 5, 5)), 1, 15) -- 4341
,( 3, E,0,0,((38,38),(29,29),( 2, 2),(99,99),(16,16),( 6, 6)), 1, 15) -- 4342
,( 3, E,0,0,((39,39),(30,30),( 3, 3),(99,99),(17,17),( 7, 7)), 1, 15) -- 4343
,( 3, E,0,0,((40,40),(31,31),( 4, 4),(99,99),(18,18),( 8, 8)), 1, 15) -- 4344
,( 3, E,0,0,((41,41),(32,32),( 5, 5),(99,99),(19,19),( 9, 9)), 1, 15) -- 4345
,( 3, E,0,0,((42,42),(33,33),( 6, 6),(99,99),(20,20),(10,10)), 1, 15) -- 4346
,( 3, E,0,0,((43,43),(34,34),( 7, 7),(99,99),(21,21),(11,11)), 1, 15) -- 4347
,( 3, E,0,0,((35,35),(27,27),( 0, 0),(99,99),(15,15),( 5, 5)), 1, 15) -- 4348
,( 3, E,0,0,((36,36),(28,28),( 1, 1),(99,99),(16,16),( 6, 6)), 1, 15) -- 4349
,( 3, E,0,0,((37,37),(29,29),( 2, 2),(99,99),(17,17),( 7, 7)), 1, 15) -- 4350
,( 3, E,0,0,((38,38),(30,30),( 3, 3),(99,99),(18,18),( 8, 8)), 1, 15) -- 4351
,( 3, E,0,0,((39,39),(31,31),( 4, 4),(99,99),(19,19),( 9, 9)), 1, 15) -- 4352
,( 3, E,0,0,((40,40),(32,32),( 5, 5),(99,99),(20,20),(10,10)), 1, 15) -- 4353
,( 3, E,0,0,((41,41),(33,33),( 6, 6),(99,99),(21,21),(11,11)), 1, 15) -- 4354
,( 3, E,0,0,((42,42),(34,34),( 7, 7),(99,99),(22,22),(12,12)), 1, 15) -- 4355
,( 3, E,0,0,((36,36),(27,27),( 0, 0),(99,99),(14,14),( 5, 5)), 1, 15) -- 4356
,( 3, E,0,0,((37,37),(28,28),( 1, 1),(99,99),(15,15),( 6, 6)), 1, 15) -- 4357
,( 3, E,0,0,((38,38),(29,29),( 2, 2),(99,99),(16,16),( 7, 7)), 1, 15) -- 4358
,( 3, E,0,0,((39,39),(30,30),( 3, 3),(99,99),(17,17),( 8, 8)), 1, 15) -- 4359
,( 3, E,0,0,((40,40),(31,31),( 4, 4),(99,99),(18,18),( 9, 9)), 1, 15) -- 4360
,( 3, E,0,0,((41,41),(32,32),( 5, 5),(99,99),(19,19),(10,10)), 1, 15) -- 4361
,( 3, E,0,0,((42,42),(33,33),( 6, 6),(99,99),(20,20),(11,11)), 1, 15) -- 4362
,( 3, E,0,0,((43,43),(34,34),( 7, 7),(99,99),(21,21),(12,12)), 1, 15) -- 4363
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(14,14),( 6, 6)), 1, 15) -- 4364
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(15,15),( 7, 7)), 1, 15) -- 4365
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(16,16),( 8, 8)), 1, 15) -- 4366
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(17,17),( 9, 9)), 1, 15) -- 4367
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(18,18),(10,10)), 1, 15) -- 4368
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(19,19),(11,11)), 1, 15) -- 4369
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(20,20),(12,12)), 1, 15) -- 4370
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(21,21),(13,13)), 1, 15) -- 4371
,( 3, E,0,0,((34,34),(25,25),( 0, 0),(99,99),(14,14),( 4, 4)), 1, 15) -- 4372
,( 3, E,0,0,((35,35),(26,26),( 1, 1),(99,99),(15,15),( 5, 5)), 1, 15) -- 4373
,( 3, E,0,0,((36,36),(27,27),( 2, 2),(99,99),(16,16),( 6, 6)), 1, 15) -- 4374
,( 3, E,0,0,((37,37),(28,28),( 3, 3),(99,99),(17,17),( 7, 7)), 1, 15) -- 4375
,( 3, E,0,0,((38,38),(29,29),( 4, 4),(99,99),(18,18),( 8, 8)), 1, 15) -- 4376
,( 3, E,0,0,((39,39),(30,30),( 5, 5),(99,99),(19,19),( 9, 9)), 1, 15) -- 4377
,( 3, E,0,0,((40,40),(31,31),( 6, 6),(99,99),(20,20),(10,10)), 1, 15) -- 4378
,( 3, E,0,0,((41,41),(32,32),( 7, 7),(99,99),(21,21),(11,11)), 1, 15) -- 4379
,( 3, E,0,0,((35,35),(26,26),( 0, 0),(99,99),(13,13),( 4, 4)), 1, 15) -- 4380
,( 3, E,0,0,((36,36),(27,27),( 1, 1),(99,99),(14,14),( 5, 5)), 1, 15) -- 4381
,( 3, E,0,0,((37,37),(28,28),( 2, 2),(99,99),(15,15),( 6, 6)), 1, 15) -- 4382
,( 3, E,0,0,((38,38),(29,29),( 3, 3),(99,99),(16,16),( 7, 7)), 1, 15) -- 4383
,( 3, E,0,0,((39,39),(30,30),( 4, 4),(99,99),(17,17),( 8, 8)), 1, 15) -- 4384
,( 3, E,0,0,((40,40),(31,31),( 5, 5),(99,99),(18,18),( 9, 9)), 1, 15) -- 4385
,( 3, E,0,0,((41,41),(32,32),( 6, 6),(99,99),(19,19),(10,10)), 1, 15) -- 4386
,( 3, E,0,0,((42,42),(33,33),( 7, 7),(99,99),(20,20),(11,11)), 1, 15) -- 4387
,( 3, E,0,0,((36,36),(27,27),( 0, 0),(99,99),(15,15),( 5, 5)), 1, 15) -- 4388
,( 3, E,0,0,((37,37),(28,28),( 1, 1),(99,99),(16,16),( 6, 6)), 1, 15) -- 4389
,( 3, E,0,0,((38,38),(29,29),( 2, 2),(99,99),(17,17),( 7, 7)), 1, 15) -- 4390
,( 3, E,0,0,((39,39),(30,30),( 3, 3),(99,99),(18,18),( 8, 8)), 1, 15) -- 4391
,( 3, E,0,0,((40,40),(31,31),( 4, 4),(99,99),(19,19),( 9, 9)), 1, 15) -- 4392
,( 3, E,0,0,((41,41),(32,32),( 5, 5),(99,99),(20,20),(10,10)), 1, 15) -- 4393
,( 3, E,0,0,((42,42),(33,33),( 6, 6),(99,99),(21,21),(11,11)), 1, 15) -- 4394
,( 3, E,0,0,((43,43),(34,34),( 7, 7),(99,99),(22,22),(12,12)), 1, 15) -- 4395
,( 3, E,0,0,((34,37),(26,27),( 0, 1),(99,99),(14,15),( 4, 7)), 1, 14) -- 4396
,( 3, E,0,0,((36,39),(28,29),( 2, 3),(99,99),(16,17),( 6, 9)), 1, 14) -- 4397
,( 3, E,0,0,((38,41),(30,31),( 4, 5),(99,99),(18,19),( 8,11)), 1, 14) -- 4398
,( 3, E,0,0,((40,43),(32,33),( 6, 7),(99,99),(20,21),(10,13)), 1, 14) -- 4399
,( 3, E,0,0,((36,39),(28,29),( 0, 1),(99,99),(14,15),( 4, 7)), 1, 14) -- 4400
,( 3, E,0,0,((38,41),(30,31),( 2, 3),(99,99),(16,17),( 6, 9)), 1, 14) -- 4401
,( 3, E,0,0,((40,43),(32,33),( 4, 5),(99,99),(18,19),( 8,11)), 1, 14) -- 4402
,( 3, E,0,0,((42,45),(34,35),( 6, 7),(99,99),(20,21),(10,13)), 1, 14) -- 4403
,( 3, E,0,0,((34,37),(26,27),( 0, 1),(99,99),(12,13),( 2, 5)), 1, 13) -- 4404
,( 3, E,0,0,((36,39),(28,29),( 2, 3),(99,99),(14,15),( 4, 7)), 1, 13) -- 4405
,( 3, E,0,0,((38,41),(30,31),( 4, 5),(99,99),(16,17),( 6, 9)), 1, 13) -- 4406
,( 3, E,0,0,((40,43),(32,33),( 6, 7),(99,99),(18,19),( 8,11)), 1, 13) -- 4407
,( 3, E,0,0,((32,35),(24,25),( 0, 1),(99,99),(14,15),( 6, 7)), 1, 13) -- 4408
,( 3, E,0,0,((34,37),(26,27),( 2, 3),(99,99),(16,17),( 8, 9)), 1, 13) -- 4409
,( 3, E,0,0,((36,39),(28,29),( 4, 5),(99,99),(18,19),(10,11)), 1, 13) -- 4410
,( 3, E,0,0,((38,41),(30,31),( 6, 7),(99,99),(20,21),(12,13)), 1, 13) -- 4411
,( 3, E,0,0,((36,39),(28,29),( 0, 1),(99,99),(12,13),( 2, 5)), 1, 12) -- 4412
,( 3, E,0,0,((38,41),(30,31),( 2, 3),(99,99),(14,15),( 4, 7)), 1, 12) -- 4413
,( 3, E,0,0,((40,43),(32,33),( 4, 5),(99,99),(16,17),( 6, 9)), 1, 12) -- 4414
,( 3, E,0,0,((42,45),(34,35),( 6, 7),(99,99),(18,19),( 8,11)), 1, 12) -- 4415
,( 3, E,0,0,((36,39),(26,27),( 0, 1),(99,99),(12,13),( 4, 7)), 1, 12) -- 4416
,( 3, E,0,0,((38,41),(28,29),( 2, 3),(99,99),(14,15),( 6, 9)), 1, 12) -- 4417
,( 3, E,0,0,((40,43),(30,31),( 4, 5),(99,99),(16,17),( 8,11)), 1, 12) -- 4418
,( 3, E,0,0,((42,45),(32,33),( 6, 7),(99,99),(18,19),(10,13)), 1, 12) -- 4419
,( 3, E,0,0,((36,39),(26,27),( 0, 1),(99,99),(14,15),( 6, 9)), 1, 12) -- 4420
,( 3, E,0,0,((38,41),(28,29),( 2, 3),(99,99),(16,17),( 8,11)), 1, 12) -- 4421
,( 3, E,0,0,((40,43),(30,31),( 4, 5),(99,99),(18,19),(10,13)), 1, 12) -- 4422
,( 3, E,0,0,((42,45),(32,33),( 6, 7),(99,99),(20,21),(12,15)), 1, 12) -- 4423
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(12,13),( 4, 7)), 1, 11) -- 4424
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(14,15),( 6, 9)), 1, 11) -- 4425
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(16,17),( 8,11)), 1, 11) -- 4426
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(18,19),(10,13)), 1, 11) -- 4427
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(14,15),( 6, 9)), 1, 11) -- 4428
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(16,17),( 8,11)), 1, 11) -- 4429
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(18,19),(10,13)), 1, 11) -- 4430
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(20,21),(12,15)), 1, 11) -- 4431
,( 3, E,0,0,((36,39),(26,27),( 0, 1),(99,99),(10,11),( 0, 3)), 1, 11) -- 4432
,( 3, E,0,0,((38,41),(28,29),( 2, 3),(99,99),(12,13),( 2, 5)), 1, 11) -- 4433
,( 3, E,0,0,((40,43),(30,31),( 4, 5),(99,99),(14,15),( 4, 7)), 1, 11) -- 4434
,( 3, E,0,0,((42,45),(32,33),( 6, 7),(99,99),(16,17),( 6, 9)), 1, 11) -- 4435
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(10,11),( 0, 3)), 1, 11) -- 4436
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(12,13),( 2, 5)), 1, 11) -- 4437
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(14,15),( 4, 7)), 1, 11) -- 4438
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(16,17),( 6, 9)), 1, 11) -- 4439
,( 3, E,0,0,((40,43),(30,31),( 0, 1),(99,99),(12,13),( 2, 5)), 1, 11) -- 4440
,( 3, E,0,0,((42,45),(32,33),( 2, 3),(99,99),(14,15),( 4, 7)), 1, 11) -- 4441
,( 3, E,0,0,((44,47),(34,35),( 4, 5),(99,99),(16,17),( 6, 9)), 1, 11) -- 4442
,( 3, E,0,0,((46,49),(36,37),( 6, 7),(99,99),(18,19),( 8,11)), 1, 11) -- 4443
,( 3, E,0,0,((38,38),(27,27),( 0, 1),(99,99),(12,13),( 2, 3)), 1, 11) -- 4444
,( 3, E,0,0,((40,40),(29,29),( 2, 3),(99,99),(14,15),( 4, 5)), 1, 11) -- 4445
,( 3, E,0,0,((42,42),(31,31),( 4, 5),(99,99),(16,17),( 6, 7)), 1, 11) -- 4446
,( 3, E,0,0,((44,44),(33,33),( 6, 7),(99,99),(18,19),( 8, 9)), 1, 11) -- 4447
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(12,13),( 0, 3)), 1, 11) -- 4448
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(14,15),( 2, 5)), 1, 11) -- 4449
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(16,17),( 4, 7)), 1, 11) -- 4450
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(18,19),( 6, 9)), 1, 11) -- 4451
,( 3, E,0,0,((40,41),(30,30),( 1, 1),(99,99),(14,14),( 4, 7)), 1, 11) -- 4452
,( 3, E,0,0,((42,43),(32,32),( 3, 3),(99,99),(16,16),( 6, 9)), 1, 11) -- 4453
,( 3, E,0,0,((44,45),(34,34),( 5, 5),(99,99),(18,18),( 8,11)), 1, 11) -- 4454
,( 3, E,0,0,((46,47),(36,36),( 7, 7),(99,99),(20,20),(10,13)), 1, 11) -- 4455
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(14,15),(10,13)), 1, 10) -- 4456
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(16,17),(12,15)), 1, 10) -- 4457
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(18,19),(14,17)), 1, 10) -- 4458
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(20,21),(16,19)), 1, 10) -- 4459
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(12,13),( 8,11)), 1, 10) -- 4460
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(14,15),(10,13)), 1, 10) -- 4461
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(16,17),(12,15)), 1, 10) -- 4462
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(18,19),(14,17)), 1, 10) -- 4463
,( 3, E,0,0,((40,43),(30,31),( 0, 1),(99,99),(12,13),( 6, 9)), 1, 10) -- 4464
,( 3, E,0,0,((42,45),(32,33),( 2, 3),(99,99),(14,15),( 8,11)), 1, 10) -- 4465
,( 3, E,0,0,((44,47),(34,35),( 4, 5),(99,99),(16,17),(10,13)), 1, 10) -- 4466
,( 3, E,0,0,((46,49),(36,37),( 6, 7),(99,99),(18,19),(12,15)), 1, 10) -- 4467
,( 3, E,0,0,((40,43),(30,31),( 1, 1),(99,99),(14,15),( 8,11)), 1, 10) -- 4468
,( 3, E,0,0,((42,45),(32,33),( 3, 3),(99,99),(16,17),(10,13)), 1, 10) -- 4469
,( 3, E,0,0,((44,47),(34,35),( 5, 5),(99,99),(18,19),(12,15)), 1, 10) -- 4470
,( 3, E,0,0,((46,49),(36,37),( 7, 7),(99,99),(20,21),(14,17)), 1, 10) -- 4471
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(10,11),( 4, 7)), 1, 10) -- 4472
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(12,13),( 6, 9)), 1, 10) -- 4473
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(14,15),( 8,11)), 1, 10) -- 4474
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(16,17),(10,13)), 1, 10) -- 4475
,( 3, E,0,0,((40,43),(30,31),( 0, 1),(99,99),(10,11),( 0, 3)), 1, 10) -- 4476
,( 3, E,0,0,((42,45),(32,33),( 2, 3),(99,99),(12,13),( 2, 5)), 1, 10) -- 4477
,( 3, E,0,0,((44,47),(34,35),( 4, 5),(99,99),(14,15),( 4, 7)), 1, 10) -- 4478
,( 3, E,0,0,((46,49),(36,37),( 6, 7),(99,99),(16,17),( 6, 9)), 1, 10) -- 4479
,( 3, E,0,0,((38,41),(28,29),( 1, 1),(99,99),(16,16),(10,13)), 1, 10) -- 4480
,( 3, E,0,0,((40,43),(30,31),( 3, 3),(99,99),(18,18),(12,15)), 1, 10) -- 4481
,( 3, E,0,0,((42,45),(32,33),( 5, 5),(99,99),(20,20),(14,17)), 1, 10) -- 4482
,( 3, E,0,0,((44,47),(34,35),( 7, 7),(99,99),(22,22),(16,19)), 1, 10) -- 4483
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),(12,13),(10,13)), 1,  9) -- 4484
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(14,15),(12,15)), 1,  9) -- 4485
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(16,17),(14,17)), 1,  9) -- 4486
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(18,19),(16,19)), 1,  9) -- 4487
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),(14,15),(12,15)), 1,  9) -- 4488
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(16,17),(14,17)), 1,  9) -- 4489
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(18,19),(16,19)), 1,  9) -- 4490
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(20,21),(18,21)), 1,  9) -- 4491
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),(10,11),( 4, 7)), 1,  9) -- 4492
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(12,13),( 6, 9)), 1,  9) -- 4493
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(14,15),( 8,11)), 1,  9) -- 4494
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(16,17),(10,13)), 1,  9) -- 4495
,( 3, E,0,0,((40,43),(28,29),( 0, 1),(99,99),(12,13),(12,15)), 1,  9) -- 4496
,( 3, E,0,0,((42,45),(30,31),( 2, 3),(99,99),(14,15),(14,17)), 1,  9) -- 4497
,( 3, E,0,0,((44,47),(32,33),( 4, 5),(99,99),(16,17),(16,19)), 1,  9) -- 4498
,( 3, E,0,0,((46,49),(34,35),( 6, 7),(99,99),(18,19),(18,21)), 1,  9) -- 4499
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(14,15),(14,17)), 1,  9) -- 4500
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(16,17),(16,19)), 1,  9) -- 4501
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(18,19),(18,21)), 1,  9) -- 4502
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(20,21),(20,23)), 1,  9) -- 4503
,( 3, E,0,0,((38,41),(28,29),( 0, 1),(99,99),(16,17),(14,17)), 1,  9) -- 4504
,( 3, E,0,0,((40,43),(30,31),( 2, 3),(99,99),(18,19),(16,19)), 1,  9) -- 4505
,( 3, E,0,0,((42,45),(32,33),( 4, 5),(99,99),(20,21),(18,21)), 1,  9) -- 4506
,( 3, E,0,0,((44,47),(34,35),( 6, 7),(99,99),(22,23),(20,23)), 1,  9) -- 4507
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),(16,17),(14,17)), 1,  9) -- 4508
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(18,19),(16,19)), 1,  9) -- 4509
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(20,21),(18,21)), 1,  9) -- 4510
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(22,23),(20,23)), 1,  9) -- 4511
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),( 8, 9),( 0, 3)), 1,  9) -- 4512
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(10,11),( 2, 5)), 1,  9) -- 4513
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(12,13),( 4, 7)), 1,  9) -- 4514
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(14,15),( 6, 9)), 1,  9) -- 4515
,( 3, E,0,0,((42,45),(30,31),( 0, 1),(99,99),(10,11),( 8,11)), 1,  9) -- 4516
,( 3, E,0,0,((44,47),(32,33),( 2, 3),(99,99),(12,13),(10,13)), 1,  9) -- 4517
,( 3, E,0,0,((46,49),(34,35),( 4, 5),(99,99),(14,15),(12,15)), 1,  9) -- 4518
,( 3, E,0,0,((48,51),(36,37),( 6, 7),(99,99),(16,17),(14,17)), 1,  9) -- 4519
,( 3, E,0,0,((40,41),(28,29),( 0, 0),(99,99),( 8, 9),( 0, 3)), 1,  9) -- 4520
,( 3, E,0,0,((42,43),(30,31),( 2, 2),(99,99),(10,11),( 2, 5)), 1,  9) -- 4521
,( 3, E,0,0,((44,45),(32,33),( 4, 4),(99,99),(12,13),( 4, 7)), 1,  9) -- 4522
,( 3, E,0,0,((46,47),(34,35),( 6, 6),(99,99),(14,15),( 6, 9)), 1,  9) -- 4523
,( 3, E,0,0,((44,45),(32,32),( 1, 1),(99,99),(10,11),( 2, 5)), 1,  9) -- 4524
,( 3, E,0,0,((46,47),(34,34),( 3, 3),(99,99),(12,13),( 4, 7)), 1,  9) -- 4525
,( 3, E,0,0,((48,49),(36,36),( 5, 5),(99,99),(14,15),( 6, 9)), 1,  9) -- 4526
,( 3, E,0,0,((50,51),(38,38),( 7, 7),(99,99),(16,17),( 8,11)), 1,  9) -- 4527
,( 3, E,0,0,((41,41),(30,30),( 1, 1),(99,99),(14,15),(12,15)), 1,  9) -- 4528
,( 3, E,0,0,((43,43),(32,32),( 3, 3),(99,99),(16,17),(14,17)), 1,  9) -- 4529
,( 3, E,0,0,((45,45),(34,34),( 5, 5),(99,99),(18,19),(16,19)), 1,  9) -- 4530
,( 3, E,0,0,((47,47),(36,36),( 7, 7),(99,99),(20,21),(18,21)), 1,  9) -- 4531
,( 3, E,0,0,((40,43),(30,31),( 0, 1),(99,99),(18,19),(18,18)), 1,  9) -- 4532
,( 3, E,0,0,((42,45),(32,33),( 2, 3),(99,99),(20,21),(20,20)), 1,  9) -- 4533
,( 3, E,0,0,((44,47),(34,35),( 4, 5),(99,99),(22,23),(22,22)), 1,  9) -- 4534
,( 3, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 8,11),(99,99)), 1,  8) -- 4535
,( 3, E,0,0,((46,49),(32,35),( 2, 3),(12,15),(10,13),(99,99)), 1,  8) -- 4536
,( 3, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(12,15),(99,99)), 1,  8) -- 4537
,( 3, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(14,17),(99,99)), 1,  8) -- 4538
,( 3, E,0,0,((44,47),(32,33),( 1, 1),(99,99),(12,15),(99,99)), 1,  8) -- 4539
,( 3, E,0,0,((46,49),(34,35),( 3, 3),(99,99),(14,17),(99,99)), 1,  8) -- 4540
,( 3, E,0,0,((48,51),(36,37),( 5, 5),(99,99),(16,19),(99,99)), 1,  8) -- 4541
,( 3, E,0,0,((50,53),(38,39),( 7, 7),(99,99),(18,21),(99,99)), 1,  8) -- 4542
,( 3, E,0,0,((44,47),(30,33),( 1, 1),(99,99),(16,19),(99,99)), 1,  8) -- 4543
,( 3, E,0,0,((46,49),(32,35),( 3, 3),(99,99),(18,21),(99,99)), 1,  8) -- 4544
,( 3, E,0,0,((48,51),(34,37),( 5, 5),(99,99),(20,23),(99,99)), 1,  8) -- 4545
,( 3, E,0,0,((50,53),(36,39),( 7, 7),(99,99),(22,25),(99,99)), 1,  8) -- 4546
,( 3, E,0,1,((42,45),(28,31),( 0, 1),(99,99),(99,99),(99,99)), 1,  7) -- 4547
,( 3, E,0,1,((44,47),(30,33),( 2, 3),(99,99),(99,99),(99,99)), 1,  7) -- 4548
,( 3, E,0,1,((46,49),(32,35),( 4, 5),(99,99),(99,99),(99,99)), 1,  7) -- 4549
,( 3, E,0,1,((48,51),(34,37),( 6, 7),(99,99),(99,99),(99,99)), 1,  7) -- 4550
,( 3, E,0,1,((44,47),(30,33),( 0, 1),(99,99),(99,99),(99,99)), 1,  7) -- 4551
,( 3, E,0,1,((46,49),(32,35),( 2, 3),(99,99),(99,99),(99,99)), 1,  7) -- 4552
,( 3, E,0,1,((48,51),(34,37),( 4, 5),(99,99),(99,99),(99,99)), 1,  7) -- 4553
,( 3, E,0,1,((50,53),(36,39),( 6, 7),(99,99),(99,99),(99,99)), 1,  7) -- 4554
,( 3, E,0,1,((54,57),(32,35),( 0, 1),(99,99),(99,99),(99,99)), 1,  7) -- 4555
,( 3, E,0,1,((56,59),(34,37),( 2, 3),(99,99),(99,99),(99,99)), 1,  7) -- 4556
,( 3, E,0,1,((58,61),(36,39),( 4, 5),(99,99),(99,99),(99,99)), 1,  7) -- 4557
,( 3, E,0,1,((60,63),(38,41),( 6, 7),(99,99),(99,99),(99,99)), 1,  7) -- 4558
,( 3, E,0,1,((38,41),(26,29),( 0, 1),(17,17),(99,99),(99,99)), 1,  6) -- 4559
,( 3, E,0,1,((40,43),(28,31),( 2, 3),(19,19),(99,99),(99,99)), 1,  6) -- 4560
,( 3, E,0,1,((42,45),(30,33),( 4, 5),(21,21),(99,99),(99,99)), 1,  6) -- 4561
,( 3, E,0,1,((44,47),(32,35),( 6, 7),(23,23),(99,99),(99,99)), 1,  6) -- 4562
,( 3, E,0,1,((42,42),(27,27),( 1, 1),(99,99),(99,99),(99,99)), 1,  5) -- 4563
,( 3, E,0,1,((44,44),(29,29),( 3, 3),(99,99),(99,99),(99,99)), 1,  5) -- 4564
,( 3, E,0,1,((46,46),(31,31),( 5, 5),(99,99),(99,99),(99,99)), 1,  5) -- 4565
,( 3, E,0,1,((48,48),(33,33),( 7, 7),(99,99),(99,99),(99,99)), 1,  5) -- 4566
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(17,17),( 8, 8)), 0, 31) -- 4567
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(18,18),( 9, 9)), 0, 31) -- 4568
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(19,19),(10,10)), 0, 31) -- 4569
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(20,20),(11,11)), 0, 31) -- 4570
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(21,21),(12,12)), 0, 31) -- 4571
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(22,22),(13,13)), 0, 31) -- 4572
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(23,23),(14,14)), 0, 31) -- 4573
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(24,24),(15,15)), 0, 31) -- 4574
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(17,17),( 8, 8)), 0, 31) -- 4575
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(18,18),( 9, 9)), 0, 31) -- 4576
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(19,19),(10,10)), 0, 31) -- 4577
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(20,20),(11,11)), 0, 31) -- 4578
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(21,21),(12,12)), 0, 31) -- 4579
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(22,22),(13,13)), 0, 31) -- 4580
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(23,23),(14,14)), 0, 31) -- 4581
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(24,24),(15,15)), 0, 31) -- 4582
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(16,16),( 8, 8)), 0, 31) -- 4583
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(17,17),( 9, 9)), 0, 31) -- 4584
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(18,18),(10,10)), 0, 31) -- 4585
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(19,19),(11,11)), 0, 31) -- 4586
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(20,20),(12,12)), 0, 31) -- 4587
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(21,21),(13,13)), 0, 31) -- 4588
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(22,22),(14,14)), 0, 31) -- 4589
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(23,23),(15,15)), 0, 31) -- 4590
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(16,16),( 7, 7)), 0, 31) -- 4591
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(17,17),( 8, 8)), 0, 31) -- 4592
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(18,18),( 9, 9)), 0, 31) -- 4593
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(19,19),(10,10)), 0, 31) -- 4594
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(20,20),(11,11)), 0, 31) -- 4595
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(21,21),(12,12)), 0, 31) -- 4596
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(22,22),(13,13)), 0, 31) -- 4597
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(23,23),(14,14)), 0, 31) -- 4598
,( 3, E,0,0,((32,32),(25,25),( 0, 0),(99,99),(17,17),( 9, 9)), 0, 31) -- 4599
,( 3, E,0,0,((33,33),(26,26),( 1, 1),(99,99),(18,18),(10,10)), 0, 31) -- 4600
,( 3, E,0,0,((34,34),(27,27),( 2, 2),(99,99),(19,19),(11,11)), 0, 31) -- 4601
,( 3, E,0,0,((35,35),(28,28),( 3, 3),(99,99),(20,20),(12,12)), 0, 31) -- 4602
,( 3, E,0,0,((36,36),(29,29),( 4, 4),(99,99),(21,21),(13,13)), 0, 31) -- 4603
,( 3, E,0,0,((37,37),(30,30),( 5, 5),(99,99),(22,22),(14,14)), 0, 31) -- 4604
,( 3, E,0,0,((38,38),(31,31),( 6, 6),(99,99),(23,23),(15,15)), 0, 31) -- 4605
,( 3, E,0,0,((39,39),(32,32),( 7, 7),(99,99),(24,24),(16,16)), 0, 31) -- 4606
,( 3, E,0,0,((32,32),(24,24),( 0, 0),(99,99),(16,16),( 8, 8)), 0, 31) -- 4607
,( 3, E,0,0,((33,33),(25,25),( 1, 1),(99,99),(17,17),( 9, 9)), 0, 31) -- 4608
,( 3, E,0,0,((34,34),(26,26),( 2, 2),(99,99),(18,18),(10,10)), 0, 31) -- 4609
,( 3, E,0,0,((35,35),(27,27),( 3, 3),(99,99),(19,19),(11,11)), 0, 31) -- 4610
,( 3, E,0,0,((36,36),(28,28),( 4, 4),(99,99),(20,20),(12,12)), 0, 31) -- 4611
,( 3, E,0,0,((37,37),(29,29),( 5, 5),(99,99),(21,21),(13,13)), 0, 31) -- 4612
,( 3, E,0,0,((38,38),(30,30),( 6, 6),(99,99),(22,22),(14,14)), 0, 31) -- 4613
,( 3, E,0,0,((39,39),(31,31),( 7, 7),(99,99),(23,23),(15,15)), 0, 31) -- 4614
,( 3, E,0,0,((32,32),(24,24),( 0, 0),(99,99),(17,17),( 8, 8)), 0, 31) -- 4615
,( 3, E,0,0,((33,33),(25,25),( 1, 1),(99,99),(18,18),( 9, 9)), 0, 31) -- 4616
,( 3, E,0,0,((34,34),(26,26),( 2, 2),(99,99),(19,19),(10,10)), 0, 31) -- 4617
,( 3, E,0,0,((35,35),(27,27),( 3, 3),(99,99),(20,20),(11,11)), 0, 31) -- 4618
,( 3, E,0,0,((36,36),(28,28),( 4, 4),(99,99),(21,21),(12,12)), 0, 31) -- 4619
,( 3, E,0,0,((37,37),(29,29),( 5, 5),(99,99),(22,22),(13,13)), 0, 31) -- 4620
,( 3, E,0,0,((38,38),(30,30),( 6, 6),(99,99),(23,23),(14,14)), 0, 31) -- 4621
,( 3, E,0,0,((39,39),(31,31),( 7, 7),(99,99),(24,24),(15,15)), 0, 31) -- 4622
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(17,17),( 9, 9)), 0, 30) -- 4623
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(18,18),(10,10)), 0, 30) -- 4624
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(19,19),(11,11)), 0, 30) -- 4625
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(20,20),(12,12)), 0, 30) -- 4626
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(21,21),(13,13)), 0, 30) -- 4627
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(22,22),(14,14)), 0, 30) -- 4628
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(23,23),(15,15)), 0, 30) -- 4629
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(24,24),(16,16)), 0, 30) -- 4630
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 24) -- 4631
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(19,19),(10,10)), 0, 24) -- 4632
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(20,20),(11,11)), 0, 24) -- 4633
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(21,21),(12,12)), 0, 24) -- 4634
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(22,22),(13,13)), 0, 24) -- 4635
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(23,23),(14,14)), 0, 24) -- 4636
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(24,24),(15,15)), 0, 24) -- 4637
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(25,25),(16,16)), 0, 24) -- 4638
,( 3, E,0,0,((30,30),(23,23),( 0, 0),(99,99),(16,16),( 8, 8)), 0, 24) -- 4639
,( 3, E,0,0,((31,31),(24,24),( 1, 1),(99,99),(17,17),( 9, 9)), 0, 24) -- 4640
,( 3, E,0,0,((32,32),(25,25),( 2, 2),(99,99),(18,18),(10,10)), 0, 24) -- 4641
,( 3, E,0,0,((33,33),(26,26),( 3, 3),(99,99),(19,19),(11,11)), 0, 24) -- 4642
,( 3, E,0,0,((34,34),(27,27),( 4, 4),(99,99),(20,20),(12,12)), 0, 24) -- 4643
,( 3, E,0,0,((35,35),(28,28),( 5, 5),(99,99),(21,21),(13,13)), 0, 24) -- 4644
,( 3, E,0,0,((36,36),(29,29),( 6, 6),(99,99),(22,22),(14,14)), 0, 24) -- 4645
,( 3, E,0,0,((37,37),(30,30),( 7, 7),(99,99),(23,23),(15,15)), 0, 24) -- 4646
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(17,17),(10,10)), 0, 24) -- 4647
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(18,18),(11,11)), 0, 24) -- 4648
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(19,19),(12,12)), 0, 24) -- 4649
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(20,20),(13,13)), 0, 24) -- 4650
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(21,21),(14,14)), 0, 24) -- 4651
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(22,22),(15,15)), 0, 24) -- 4652
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(23,23),(16,16)), 0, 24) -- 4653
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(24,24),(17,17)), 0, 24) -- 4654
,( 3, E,0,0,((30,30),(24,24),( 0, 0),(99,99),(17,17),( 8, 8)), 0, 23) -- 4655
,( 3, E,0,0,((31,31),(25,25),( 1, 1),(99,99),(18,18),( 9, 9)), 0, 23) -- 4656
,( 3, E,0,0,((32,32),(26,26),( 2, 2),(99,99),(19,19),(10,10)), 0, 23) -- 4657
,( 3, E,0,0,((33,33),(27,27),( 3, 3),(99,99),(20,20),(11,11)), 0, 23) -- 4658
,( 3, E,0,0,((34,34),(28,28),( 4, 4),(99,99),(21,21),(12,12)), 0, 23) -- 4659
,( 3, E,0,0,((35,35),(29,29),( 5, 5),(99,99),(22,22),(13,13)), 0, 23) -- 4660
,( 3, E,0,0,((36,36),(30,30),( 6, 6),(99,99),(23,23),(14,14)), 0, 23) -- 4661
,( 3, E,0,0,((37,37),(31,31),( 7, 7),(99,99),(24,24),(15,15)), 0, 23) -- 4662
,( 3, E,0,0,((30,30),(23,23),( 0, 0),(99,99),(17,17),( 8, 8)), 0, 23) -- 4663
,( 3, E,0,0,((31,31),(24,24),( 1, 1),(99,99),(18,18),( 9, 9)), 0, 23) -- 4664
,( 3, E,0,0,((32,32),(25,25),( 2, 2),(99,99),(19,19),(10,10)), 0, 23) -- 4665
,( 3, E,0,0,((33,33),(26,26),( 3, 3),(99,99),(20,20),(11,11)), 0, 23) -- 4666
,( 3, E,0,0,((34,34),(27,27),( 4, 4),(99,99),(21,21),(12,12)), 0, 23) -- 4667
,( 3, E,0,0,((35,35),(28,28),( 5, 5),(99,99),(22,22),(13,13)), 0, 23) -- 4668
,( 3, E,0,0,((36,36),(29,29),( 6, 6),(99,99),(23,23),(14,14)), 0, 23) -- 4669
,( 3, E,0,0,((37,37),(30,30),( 7, 7),(99,99),(24,24),(15,15)), 0, 23) -- 4670
,( 3, E,0,0,((30,30),(24,24),( 0, 0),(99,99),(17,17),( 9, 9)), 0, 22) -- 4671
,( 3, E,0,0,((31,31),(25,25),( 1, 1),(99,99),(18,18),(10,10)), 0, 22) -- 4672
,( 3, E,0,0,((32,32),(26,26),( 2, 2),(99,99),(19,19),(11,11)), 0, 22) -- 4673
,( 3, E,0,0,((33,33),(27,27),( 3, 3),(99,99),(20,20),(12,12)), 0, 22) -- 4674
,( 3, E,0,0,((34,34),(28,28),( 4, 4),(99,99),(21,21),(13,13)), 0, 22) -- 4675
,( 3, E,0,0,((35,35),(29,29),( 5, 5),(99,99),(22,22),(14,14)), 0, 22) -- 4676
,( 3, E,0,0,((36,36),(30,30),( 6, 6),(99,99),(23,23),(15,15)), 0, 22) -- 4677
,( 3, E,0,0,((37,37),(31,31),( 7, 7),(99,99),(24,24),(16,16)), 0, 22) -- 4678
,( 3, E,0,0,((30,30),(23,23),( 0, 0),(99,99),(17,17),( 9, 9)), 0, 22) -- 4679
,( 3, E,0,0,((31,31),(24,24),( 1, 1),(99,99),(18,18),(10,10)), 0, 22) -- 4680
,( 3, E,0,0,((32,32),(25,25),( 2, 2),(99,99),(19,19),(11,11)), 0, 22) -- 4681
,( 3, E,0,0,((33,33),(26,26),( 3, 3),(99,99),(20,20),(12,12)), 0, 22) -- 4682
,( 3, E,0,0,((34,34),(27,27),( 4, 4),(99,99),(21,21),(13,13)), 0, 22) -- 4683
,( 3, E,0,0,((35,35),(28,28),( 5, 5),(99,99),(22,22),(14,14)), 0, 22) -- 4684
,( 3, E,0,0,((36,36),(29,29),( 6, 6),(99,99),(23,23),(15,15)), 0, 22) -- 4685
,( 3, E,0,0,((37,37),(30,30),( 7, 7),(99,99),(24,24),(16,16)), 0, 22) -- 4686
,( 3, E,0,0,((30,30),(24,24),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 20) -- 4687
,( 3, E,0,0,((31,31),(25,25),( 1, 1),(99,99),(19,19),(10,10)), 0, 20) -- 4688
,( 3, E,0,0,((32,32),(26,26),( 2, 2),(99,99),(20,20),(11,11)), 0, 20) -- 4689
,( 3, E,0,0,((33,33),(27,27),( 3, 3),(99,99),(21,21),(12,12)), 0, 20) -- 4690
,( 3, E,0,0,((34,34),(28,28),( 4, 4),(99,99),(22,22),(13,13)), 0, 20) -- 4691
,( 3, E,0,0,((35,35),(29,29),( 5, 5),(99,99),(23,23),(14,14)), 0, 20) -- 4692
,( 3, E,0,0,((36,36),(30,30),( 6, 6),(99,99),(24,24),(15,15)), 0, 20) -- 4693
,( 3, E,0,0,((37,37),(31,31),( 7, 7),(99,99),(25,25),(16,16)), 0, 20) -- 4694
,( 3, E,0,0,((31,31),(24,24),( 0, 0),(99,99),(18,18),(10,10)), 0, 20) -- 4695
,( 3, E,0,0,((32,32),(25,25),( 1, 1),(99,99),(19,19),(11,11)), 0, 20) -- 4696
,( 3, E,0,0,((33,33),(26,26),( 2, 2),(99,99),(20,20),(12,12)), 0, 20) -- 4697
,( 3, E,0,0,((34,34),(27,27),( 3, 3),(99,99),(21,21),(13,13)), 0, 20) -- 4698
,( 3, E,0,0,((35,35),(28,28),( 4, 4),(99,99),(22,22),(14,14)), 0, 20) -- 4699
,( 3, E,0,0,((36,36),(29,29),( 5, 5),(99,99),(23,23),(15,15)), 0, 20) -- 4700
,( 3, E,0,0,((37,37),(30,30),( 6, 6),(99,99),(24,24),(16,16)), 0, 20) -- 4701
,( 3, E,0,0,((38,38),(31,31),( 7, 7),(99,99),(25,25),(17,17)), 0, 20) -- 4702
,( 3, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 4703
,( 3, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 4704
,( 3, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 4705
,( 3, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 4706
,( 3, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 4707
,( 3, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 4708
,( 3, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 4709
,( 3, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 4710
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 18) -- 4711
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 18) -- 4712
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 18) -- 4713
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 18) -- 4714
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 18) -- 4715
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 18) -- 4716
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 18) -- 4717
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 18) -- 4718
,( 3, E,0,0,((30,30),(23,23),( 0, 0),(99,99),(18,18),(10,10)), 0, 18) -- 4719
,( 3, E,0,0,((31,31),(24,24),( 1, 1),(99,99),(19,19),(11,11)), 0, 18) -- 4720
,( 3, E,0,0,((32,32),(25,25),( 2, 2),(99,99),(20,20),(12,12)), 0, 18) -- 4721
,( 3, E,0,0,((33,33),(26,26),( 3, 3),(99,99),(21,21),(13,13)), 0, 18) -- 4722
,( 3, E,0,0,((34,34),(27,27),( 4, 4),(99,99),(22,22),(14,14)), 0, 18) -- 4723
,( 3, E,0,0,((35,35),(28,28),( 5, 5),(99,99),(23,23),(15,15)), 0, 18) -- 4724
,( 3, E,0,0,((36,36),(29,29),( 6, 6),(99,99),(24,24),(16,16)), 0, 18) -- 4725
,( 3, E,0,0,((37,37),(30,30),( 7, 7),(99,99),(25,25),(17,17)), 0, 18) -- 4726
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 18) -- 4727
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(99,99),(19,19),(10,10)), 0, 18) -- 4728
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(99,99),(20,20),(11,11)), 0, 18) -- 4729
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(99,99),(21,21),(12,12)), 0, 18) -- 4730
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(99,99),(22,22),(13,13)), 0, 18) -- 4731
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(99,99),(23,23),(14,14)), 0, 18) -- 4732
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(99,99),(24,24),(15,15)), 0, 18) -- 4733
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(99,99),(25,25),(16,16)), 0, 18) -- 4734
,( 3, E,0,0,((30,30),(23,23),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 18) -- 4735
,( 3, E,0,0,((31,31),(24,24),( 1, 1),(99,99),(19,19),(10,10)), 0, 18) -- 4736
,( 3, E,0,0,((32,32),(25,25),( 2, 2),(99,99),(20,20),(11,11)), 0, 18) -- 4737
,( 3, E,0,0,((33,33),(26,26),( 3, 3),(99,99),(21,21),(12,12)), 0, 18) -- 4738
,( 3, E,0,0,((34,34),(27,27),( 4, 4),(99,99),(22,22),(13,13)), 0, 18) -- 4739
,( 3, E,0,0,((35,35),(28,28),( 5, 5),(99,99),(23,23),(14,14)), 0, 18) -- 4740
,( 3, E,0,0,((36,36),(29,29),( 6, 6),(99,99),(24,24),(15,15)), 0, 18) -- 4741
,( 3, E,0,0,((37,37),(30,30),( 7, 7),(99,99),(25,25),(16,16)), 0, 18) -- 4742
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(99,99),(17,17),( 9, 9)), 0, 18) -- 4743
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(99,99),(18,18),(10,10)), 0, 18) -- 4744
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(99,99),(19,19),(11,11)), 0, 18) -- 4745
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(99,99),(20,20),(12,12)), 0, 18) -- 4746
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(99,99),(21,21),(13,13)), 0, 18) -- 4747
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(99,99),(22,22),(14,14)), 0, 18) -- 4748
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(99,99),(23,23),(15,15)), 0, 18) -- 4749
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(99,99),(24,24),(16,16)), 0, 18) -- 4750
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(99,99),(19,19),(11,11)), 0, 17) -- 4751
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(99,99),(20,20),(12,12)), 0, 17) -- 4752
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(99,99),(21,21),(13,13)), 0, 17) -- 4753
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(99,99),(22,22),(14,14)), 0, 17) -- 4754
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(99,99),(23,23),(15,15)), 0, 17) -- 4755
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(99,99),(24,24),(16,16)), 0, 17) -- 4756
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(99,99),(25,25),(17,17)), 0, 17) -- 4757
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(99,99),(26,26),(18,18)), 0, 17) -- 4758
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(99,99),(18,18),(11,11)), 0, 17) -- 4759
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(99,99),(19,19),(12,12)), 0, 17) -- 4760
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(99,99),(20,20),(13,13)), 0, 17) -- 4761
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(99,99),(21,21),(14,14)), 0, 17) -- 4762
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(99,99),(22,22),(15,15)), 0, 17) -- 4763
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(99,99),(23,23),(16,16)), 0, 17) -- 4764
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(99,99),(24,24),(17,17)), 0, 17) -- 4765
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(99,99),(25,25),(18,18)), 0, 17) -- 4766
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(99,99),(19,19),(10,10)), 0, 17) -- 4767
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(99,99),(20,20),(11,11)), 0, 17) -- 4768
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(99,99),(21,21),(12,12)), 0, 17) -- 4769
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(99,99),(22,22),(13,13)), 0, 17) -- 4770
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(99,99),(23,23),(14,14)), 0, 17) -- 4771
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(99,99),(24,24),(15,15)), 0, 17) -- 4772
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(99,99),(25,25),(16,16)), 0, 17) -- 4773
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(99,99),(26,26),(17,17)), 0, 17) -- 4774
,( 3, E,0,0,((30,30),(24,24),( 0, 0),(99,99),(19,19),(10,10)), 0, 17) -- 4775
,( 3, E,0,0,((31,31),(25,25),( 1, 1),(99,99),(20,20),(11,11)), 0, 17) -- 4776
,( 3, E,0,0,((32,32),(26,26),( 2, 2),(99,99),(21,21),(12,12)), 0, 17) -- 4777
,( 3, E,0,0,((33,33),(27,27),( 3, 3),(99,99),(22,22),(13,13)), 0, 17) -- 4778
,( 3, E,0,0,((34,34),(28,28),( 4, 4),(99,99),(23,23),(14,14)), 0, 17) -- 4779
,( 3, E,0,0,((35,35),(29,29),( 5, 5),(99,99),(24,24),(15,15)), 0, 17) -- 4780
,( 3, E,0,0,((36,36),(30,30),( 6, 6),(99,99),(25,25),(16,16)), 0, 17) -- 4781
,( 3, E,0,0,((37,37),(31,31),( 7, 7),(99,99),(26,26),(17,17)), 0, 17) -- 4782
,( 3, E,0,0,((29,29),(22,22),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 17) -- 4783
,( 3, E,0,0,((30,30),(23,23),( 1, 1),(99,99),(19,19),(10,10)), 0, 17) -- 4784
,( 3, E,0,0,((31,31),(24,24),( 2, 2),(99,99),(20,20),(11,11)), 0, 17) -- 4785
,( 3, E,0,0,((32,32),(25,25),( 3, 3),(99,99),(21,21),(12,12)), 0, 17) -- 4786
,( 3, E,0,0,((33,33),(26,26),( 4, 4),(99,99),(22,22),(13,13)), 0, 17) -- 4787
,( 3, E,0,0,((34,34),(27,27),( 5, 5),(99,99),(23,23),(14,14)), 0, 17) -- 4788
,( 3, E,0,0,((35,35),(28,28),( 6, 6),(99,99),(24,24),(15,15)), 0, 17) -- 4789
,( 3, E,0,0,((36,36),(29,29),( 7, 7),(99,99),(25,25),(16,16)), 0, 17) -- 4790
,( 3, E,0,0,((28,28),(22,22),( 0, 0),(99,99),(18,18),(11,11)), 0, 16) -- 4791
,( 3, E,0,0,((29,29),(23,23),( 1, 1),(99,99),(19,19),(12,12)), 0, 16) -- 4792
,( 3, E,0,0,((30,30),(24,24),( 2, 2),(99,99),(20,20),(13,13)), 0, 16) -- 4793
,( 3, E,0,0,((31,31),(25,25),( 3, 3),(99,99),(21,21),(14,14)), 0, 16) -- 4794
,( 3, E,0,0,((32,32),(26,26),( 4, 4),(99,99),(22,22),(15,15)), 0, 16) -- 4795
,( 3, E,0,0,((33,33),(27,27),( 5, 5),(99,99),(23,23),(16,16)), 0, 16) -- 4796
,( 3, E,0,0,((34,34),(28,28),( 6, 6),(99,99),(24,24),(17,17)), 0, 16) -- 4797
,( 3, E,0,0,((35,35),(29,29),( 7, 7),(99,99),(25,25),(18,18)), 0, 16) -- 4798
,( 3, E,0,0,((28,28),(23,23),( 0, 0),(99,99),(18,18),(10,10)), 0, 16) -- 4799
,( 3, E,0,0,((29,29),(24,24),( 1, 1),(99,99),(19,19),(11,11)), 0, 16) -- 4800
,( 3, E,0,0,((30,30),(25,25),( 2, 2),(99,99),(20,20),(12,12)), 0, 16) -- 4801
,( 3, E,0,0,((31,31),(26,26),( 3, 3),(99,99),(21,21),(13,13)), 0, 16) -- 4802
,( 3, E,0,0,((32,32),(27,27),( 4, 4),(99,99),(22,22),(14,14)), 0, 16) -- 4803
,( 3, E,0,0,((33,33),(28,28),( 5, 5),(99,99),(23,23),(15,15)), 0, 16) -- 4804
,( 3, E,0,0,((34,34),(29,29),( 6, 6),(99,99),(24,24),(16,16)), 0, 16) -- 4805
,( 3, E,0,0,((35,35),(30,30),( 7, 7),(99,99),(25,25),(17,17)), 0, 16) -- 4806
,( 3, E,0,0,((28,28),(23,23),( 0, 0),(99,99),(19,19),(11,11)), 0, 16) -- 4807
,( 3, E,0,0,((29,29),(24,24),( 1, 1),(99,99),(20,20),(12,12)), 0, 16) -- 4808
,( 3, E,0,0,((30,30),(25,25),( 2, 2),(99,99),(21,21),(13,13)), 0, 16) -- 4809
,( 3, E,0,0,((31,31),(26,26),( 3, 3),(99,99),(22,22),(14,14)), 0, 16) -- 4810
,( 3, E,0,0,((32,32),(27,27),( 4, 4),(99,99),(23,23),(15,15)), 0, 16) -- 4811
,( 3, E,0,0,((33,33),(28,28),( 5, 5),(99,99),(24,24),(16,16)), 0, 16) -- 4812
,( 3, E,0,0,((34,34),(29,29),( 6, 6),(99,99),(25,25),(17,17)), 0, 16) -- 4813
,( 3, E,0,0,((35,35),(30,30),( 7, 7),(99,99),(26,26),(18,18)), 0, 16) -- 4814
,( 3, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(99,99),(11,11)), 0, 16) -- 4815
,( 3, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(99,99),(12,12)), 0, 16) -- 4816
,( 3, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(99,99),(13,13)), 0, 16) -- 4817
,( 3, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(99,99),(14,14)), 0, 16) -- 4818
,( 3, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(99,99),(15,15)), 0, 16) -- 4819
,( 3, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(99,99),(16,16)), 0, 16) -- 4820
,( 3, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(99,99),(17,17)), 0, 16) -- 4821
,( 3, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(99,99),(18,18)), 0, 16) -- 4822
,( 3, E,0,0,((28,28),(23,23),( 0, 0),(99,99),(19,19),(10,10)), 0, 15) -- 4823
,( 3, E,0,0,((29,29),(24,24),( 1, 1),(99,99),(20,20),(11,11)), 0, 15) -- 4824
,( 3, E,0,0,((30,30),(25,25),( 2, 2),(99,99),(21,21),(12,12)), 0, 15) -- 4825
,( 3, E,0,0,((31,31),(26,26),( 3, 3),(99,99),(22,22),(13,13)), 0, 15) -- 4826
,( 3, E,0,0,((32,32),(27,27),( 4, 4),(99,99),(23,23),(14,14)), 0, 15) -- 4827
,( 3, E,0,0,((33,33),(28,28),( 5, 5),(99,99),(24,24),(15,15)), 0, 15) -- 4828
,( 3, E,0,0,((34,34),(29,29),( 6, 6),(99,99),(25,25),(16,16)), 0, 15) -- 4829
,( 3, E,0,0,((35,35),(30,30),( 7, 7),(99,99),(26,26),(17,17)), 0, 15) -- 4830
,( 3, E,0,0,((28,28),(22,22),( 0, 0),(99,99),(19,19),(11,11)), 0, 15) -- 4831
,( 3, E,0,0,((29,29),(23,23),( 1, 1),(99,99),(20,20),(12,12)), 0, 15) -- 4832
,( 3, E,0,0,((30,30),(24,24),( 2, 2),(99,99),(21,21),(13,13)), 0, 15) -- 4833
,( 3, E,0,0,((31,31),(25,25),( 3, 3),(99,99),(22,22),(14,14)), 0, 15) -- 4834
,( 3, E,0,0,((32,32),(26,26),( 4, 4),(99,99),(23,23),(15,15)), 0, 15) -- 4835
,( 3, E,0,0,((33,33),(27,27),( 5, 5),(99,99),(24,24),(16,16)), 0, 15) -- 4836
,( 3, E,0,0,((34,34),(28,28),( 6, 6),(99,99),(25,25),(17,17)), 0, 15) -- 4837
,( 3, E,0,0,((35,35),(29,29),( 7, 7),(99,99),(26,26),(18,18)), 0, 15) -- 4838
,( 3, E,0,0,((28,28),(23,23),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 15) -- 4839
,( 3, E,0,0,((29,29),(24,24),( 1, 1),(99,99),(19,19),(10,10)), 0, 15) -- 4840
,( 3, E,0,0,((30,30),(25,25),( 2, 2),(99,99),(20,20),(11,11)), 0, 15) -- 4841
,( 3, E,0,0,((31,31),(26,26),( 3, 3),(99,99),(21,21),(12,12)), 0, 15) -- 4842
,( 3, E,0,0,((32,32),(27,27),( 4, 4),(99,99),(22,22),(13,13)), 0, 15) -- 4843
,( 3, E,0,0,((33,33),(28,28),( 5, 5),(99,99),(23,23),(14,14)), 0, 15) -- 4844
,( 3, E,0,0,((34,34),(29,29),( 6, 6),(99,99),(24,24),(15,15)), 0, 15) -- 4845
,( 3, E,0,0,((35,35),(30,30),( 7, 7),(99,99),(25,25),(16,16)), 0, 15) -- 4846
,( 3, E,0,0,((28,28),(22,22),( 0, 0),(99,99),(18,18),(10,10)), 0, 15) -- 4847
,( 3, E,0,0,((29,29),(23,23),( 1, 1),(99,99),(19,19),(11,11)), 0, 15) -- 4848
,( 3, E,0,0,((30,30),(24,24),( 2, 2),(99,99),(20,20),(12,12)), 0, 15) -- 4849
,( 3, E,0,0,((31,31),(25,25),( 3, 3),(99,99),(21,21),(13,13)), 0, 15) -- 4850
,( 3, E,0,0,((32,32),(26,26),( 4, 4),(99,99),(22,22),(14,14)), 0, 15) -- 4851
,( 3, E,0,0,((33,33),(27,27),( 5, 5),(99,99),(23,23),(15,15)), 0, 15) -- 4852
,( 3, E,0,0,((34,34),(28,28),( 6, 6),(99,99),(24,24),(16,16)), 0, 15) -- 4853
,( 3, E,0,0,((35,35),(29,29),( 7, 7),(99,99),(25,25),(17,17)), 0, 15) -- 4854
,( 3, E,0,0,((28,28),(22,22),( 0, 0),(99,99),(18,18),( 9, 9)), 0, 15) -- 4855
,( 3, E,0,0,((29,29),(23,23),( 1, 1),(99,99),(19,19),(10,10)), 0, 15) -- 4856
,( 3, E,0,0,((30,30),(24,24),( 2, 2),(99,99),(20,20),(11,11)), 0, 15) -- 4857
,( 3, E,0,0,((31,31),(25,25),( 3, 3),(99,99),(21,21),(12,12)), 0, 15) -- 4858
,( 3, E,0,0,((32,32),(26,26),( 4, 4),(99,99),(22,22),(13,13)), 0, 15) -- 4859
,( 3, E,0,0,((33,33),(27,27),( 5, 5),(99,99),(23,23),(14,14)), 0, 15) -- 4860
,( 3, E,0,0,((34,34),(28,28),( 6, 6),(99,99),(24,24),(15,15)), 0, 15) -- 4861
,( 3, E,0,0,((35,35),(29,29),( 7, 7),(99,99),(25,25),(16,16)), 0, 15) -- 4862
,( 3, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(18,19),(10,13)), 0, 14) -- 4863
,( 3, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(20,21),(12,15)), 0, 14) -- 4864
,( 3, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(22,23),(14,17)), 0, 14) -- 4865
,( 3, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(24,25),(16,19)), 0, 14) -- 4866
,( 3, E,0,0,((26,29),(22,23),( 0, 1),(99,99),(20,21),(10,13)), 0, 14) -- 4867
,( 3, E,0,0,((28,31),(24,25),( 2, 3),(99,99),(22,23),(12,15)), 0, 14) -- 4868
,( 3, E,0,0,((30,33),(26,27),( 4, 5),(99,99),(24,25),(14,17)), 0, 14) -- 4869
,( 3, E,0,0,((32,35),(28,29),( 6, 7),(99,99),(26,27),(16,19)), 0, 14) -- 4870
,( 3, E,0,0,((28,31),(24,24),( 1, 1),(99,99),(20,21),(10,13)), 0, 14) -- 4871
,( 3, E,0,0,((30,33),(26,26),( 3, 3),(99,99),(22,23),(12,15)), 0, 14) -- 4872
,( 3, E,0,0,((32,35),(28,28),( 5, 5),(99,99),(24,25),(14,17)), 0, 14) -- 4873
,( 3, E,0,0,((34,37),(30,30),( 7, 7),(99,99),(26,27),(16,19)), 0, 14) -- 4874
,( 3, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(18,19),( 8, 9)), 0, 13) -- 4875
,( 3, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(20,21),(10,11)), 0, 13) -- 4876
,( 3, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(22,23),(12,13)), 0, 13) -- 4877
,( 3, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(24,25),(14,15)), 0, 13) -- 4878
,( 3, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(99,99),(10,13)), 0, 13) -- 4879
,( 3, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(99,99),(12,15)), 0, 13) -- 4880
,( 3, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(99,99),(14,17)), 0, 13) -- 4881
,( 3, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(99,99),(16,19)), 0, 13) -- 4882
,( 3, E,0,0,((24,27),(21,21),( 0, 0),(99,99),(19,19),(10,13)), 0, 13) -- 4883
,( 3, E,0,0,((26,29),(23,23),( 2, 2),(99,99),(21,21),(12,15)), 0, 13) -- 4884
,( 3, E,0,0,((28,31),(25,25),( 4, 4),(99,99),(23,23),(14,17)), 0, 13) -- 4885
,( 3, E,0,0,((30,33),(27,27),( 6, 6),(99,99),(25,25),(16,19)), 0, 13) -- 4886
,( 3, E,0,0,((28,31),(24,24),( 1, 1),(99,99),(22,22),(12,15)), 0, 13) -- 4887
,( 3, E,0,0,((30,33),(26,26),( 3, 3),(99,99),(24,24),(14,17)), 0, 13) -- 4888
,( 3, E,0,0,((32,35),(28,28),( 5, 5),(99,99),(26,26),(16,19)), 0, 13) -- 4889
,( 3, E,0,0,((34,37),(30,30),( 7, 7),(99,99),(28,28),(18,21)), 0, 13) -- 4890
,( 3, E,0,0,((24,27),(20,21),( 0, 1),(99,99),(20,21),(10,13)), 0, 12) -- 4891
,( 3, E,0,0,((26,29),(22,23),( 2, 3),(99,99),(22,23),(12,15)), 0, 12) -- 4892
,( 3, E,0,0,((28,31),(24,25),( 4, 5),(99,99),(24,25),(14,17)), 0, 12) -- 4893
,( 3, E,0,0,((30,33),(26,27),( 6, 7),(99,99),(26,27),(16,19)), 0, 12) -- 4894
,( 3, E,0,0,((26,29),(22,23),( 1, 1),(99,99),(22,23),(12,15)), 0, 12) -- 4895
,( 3, E,0,0,((28,31),(24,25),( 3, 3),(99,99),(24,25),(14,17)), 0, 12) -- 4896
,( 3, E,0,0,((30,33),(26,27),( 5, 5),(99,99),(26,27),(16,19)), 0, 12) -- 4897
,( 3, E,0,0,((32,35),(28,29),( 7, 7),(99,99),(28,29),(18,21)), 0, 12) -- 4898
,( 3, E,0,0,((24,27),(21,21),( 0, 0),(17,17),(99,99),(10,13)), 0, 12) -- 4899
,( 3, E,0,0,((26,29),(23,23),( 2, 2),(19,19),(99,99),(12,15)), 0, 12) -- 4900
,( 3, E,0,0,((28,31),(25,25),( 4, 4),(21,21),(99,99),(14,17)), 0, 12) -- 4901
,( 3, E,0,0,((30,33),(27,27),( 6, 6),(23,23),(99,99),(16,19)), 0, 12) -- 4902
,( 3, E,0,0,((26,29),(22,23),( 0, 1),(99,99),(21,21),(14,15)), 0, 12) -- 4903
,( 3, E,0,0,((28,31),(24,25),( 2, 3),(99,99),(23,23),(16,17)), 0, 12) -- 4904
,( 3, E,0,0,((30,33),(26,27),( 4, 5),(99,99),(25,25),(18,19)), 0, 12) -- 4905
,( 3, E,0,0,((32,35),(28,29),( 6, 7),(99,99),(27,27),(20,21)), 0, 12) -- 4906
,( 3, E,0,0,((24,27),(22,23),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 4907
,( 3, E,0,0,((26,29),(24,25),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 4908
,( 3, E,0,0,((28,31),(26,27),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 4909
,( 3, E,0,0,((30,33),(28,29),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 4910
,( 3, E,0,0,((24,27),(20,21),( 0, 1),(18,18),(18,19),( 6, 9)), 0, 11) -- 4911
,( 3, E,0,0,((26,29),(22,23),( 2, 3),(20,20),(20,21),( 8,11)), 0, 11) -- 4912
,( 3, E,0,0,((28,31),(24,25),( 4, 5),(22,22),(22,23),(10,13)), 0, 11) -- 4913
,( 3, E,0,0,((30,33),(26,27),( 6, 7),(24,24),(24,25),(12,15)), 0, 11) -- 4914
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(99,99),(10,13)), 0, 11) -- 4915
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(99,99),(12,15)), 0, 11) -- 4916
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(99,99),(14,17)), 0, 11) -- 4917
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(99,99),(16,19)), 0, 11) -- 4918
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(22,23),(12,15)), 0, 11) -- 4919
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(24,25),(14,17)), 0, 11) -- 4920
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(26,27),(16,19)), 0, 11) -- 4921
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(28,29),(18,21)), 0, 11) -- 4922
,( 3, E,0,0,((25,25),(22,22),( 0, 1),(99,99),(22,23),(12,15)), 0, 11) -- 4923
,( 3, E,0,0,((27,27),(24,24),( 2, 3),(99,99),(24,25),(14,17)), 0, 11) -- 4924
,( 3, E,0,0,((29,29),(26,26),( 4, 5),(99,99),(26,27),(16,19)), 0, 11) -- 4925
,( 3, E,0,0,((31,31),(28,28),( 6, 7),(99,99),(28,29),(18,21)), 0, 11) -- 4926
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(20,21),( 6, 9)), 0, 11) -- 4927
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(22,23),( 8,11)), 0, 11) -- 4928
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(24,25),(10,13)), 0, 11) -- 4929
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(26,27),(12,15)), 0, 11) -- 4930
,( 3, E,0,0,((24,27),(22,22),( 1, 1),(18,19),(99,99),(12,15)), 0, 11) -- 4931
,( 3, E,0,0,((26,29),(24,24),( 3, 3),(20,21),(99,99),(14,17)), 0, 11) -- 4932
,( 3, E,0,0,((28,31),(26,26),( 5, 5),(22,23),(99,99),(16,19)), 0, 11) -- 4933
,( 3, E,0,0,((30,33),(28,28),( 7, 7),(24,25),(99,99),(18,21)), 0, 11) -- 4934
,( 3, E,0,0,((24,27),(22,23),( 1, 1),(99,99),(24,24),(14,17)), 0, 11) -- 4935
,( 3, E,0,0,((26,29),(24,25),( 3, 3),(99,99),(26,26),(16,19)), 0, 11) -- 4936
,( 3, E,0,0,((28,31),(26,27),( 5, 5),(99,99),(28,28),(18,21)), 0, 11) -- 4937
,( 3, E,0,0,((30,33),(28,29),( 7, 7),(99,99),(30,30),(20,23)), 0, 11) -- 4938
,( 3, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(99,99),( 8,11)), 0, 11) -- 4939
,( 3, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(99,99),(10,13)), 0, 11) -- 4940
,( 3, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(99,99),(12,15)), 0, 11) -- 4941
,( 3, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(99,99),(14,17)), 0, 11) -- 4942
,( 3, E,0,0,((25,25),(22,22),( 0, 1),(99,99),(21,21),(12,15)), 0, 11) -- 4943
,( 3, E,0,0,((27,27),(24,24),( 2, 3),(99,99),(23,23),(14,17)), 0, 11) -- 4944
,( 3, E,0,0,((29,29),(26,26),( 4, 5),(99,99),(25,25),(16,19)), 0, 11) -- 4945
,( 3, E,0,0,((31,31),(28,28),( 6, 7),(99,99),(27,27),(18,21)), 0, 11) -- 4946
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 4, 7)), 0, 10) -- 4947
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 6, 9)), 0, 10) -- 4948
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 8,11)), 0, 10) -- 4949
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),(10,13)), 0, 10) -- 4950
,( 3, E,0,0,((20,23),(18,19),( 0, 1),(99,99),(20,21),( 8,11)), 0, 10) -- 4951
,( 3, E,0,0,((22,25),(20,21),( 2, 3),(99,99),(22,23),(10,13)), 0, 10) -- 4952
,( 3, E,0,0,((24,27),(22,23),( 4, 5),(99,99),(24,25),(12,15)), 0, 10) -- 4953
,( 3, E,0,0,((26,29),(24,25),( 6, 7),(99,99),(26,27),(14,17)), 0, 10) -- 4954
,( 3, E,0,0,((24,27),(22,22),( 1, 1),(99,99),(22,23),( 8,11)), 0, 10) -- 4955
,( 3, E,0,0,((26,29),(24,24),( 3, 3),(99,99),(24,25),(10,13)), 0, 10) -- 4956
,( 3, E,0,0,((28,31),(26,26),( 5, 5),(99,99),(26,27),(12,15)), 0, 10) -- 4957
,( 3, E,0,0,((30,33),(28,28),( 7, 7),(99,99),(28,29),(14,17)), 0, 10) -- 4958
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(99,99),( 8, 9)), 0, 10) -- 4959
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(99,99),(10,11)), 0, 10) -- 4960
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(99,99),(12,13)), 0, 10) -- 4961
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(99,99),(14,15)), 0, 10) -- 4962
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(22,23),( 8,11)), 0, 10) -- 4963
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(24,25),(10,13)), 0, 10) -- 4964
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(26,27),(12,15)), 0, 10) -- 4965
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(28,29),(14,17)), 0, 10) -- 4966
,( 3, E,0,0,((22,23),(20,21),( 0, 1),(99,99),(20,21),(10,13)), 0, 10) -- 4967
,( 3, E,0,0,((24,25),(22,23),( 2, 3),(99,99),(22,23),(12,15)), 0, 10) -- 4968
,( 3, E,0,0,((26,27),(24,25),( 4, 5),(99,99),(24,25),(14,17)), 0, 10) -- 4969
,( 3, E,0,0,((28,29),(26,27),( 6, 7),(99,99),(26,27),(16,19)), 0, 10) -- 4970
,( 3, E,0,0,((24,27),(22,23),( 0, 1),(99,99),(18,19),( 4, 7)), 0, 10) -- 4971
,( 3, E,0,0,((26,29),(24,25),( 2, 3),(99,99),(20,21),( 6, 9)), 0, 10) -- 4972
,( 3, E,0,0,((28,31),(26,27),( 4, 5),(99,99),(22,23),( 8,11)), 0, 10) -- 4973
,( 3, E,0,0,((30,33),(28,29),( 6, 7),(99,99),(24,25),(10,13)), 0, 10) -- 4974
,( 3, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(99,99),(10,13)), 0, 10) -- 4975
,( 3, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(99,99),(12,15)), 0, 10) -- 4976
,( 3, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(99,99),(14,17)), 0, 10) -- 4977
,( 3, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(99,99),(16,19)), 0, 10) -- 4978
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(16,17),( 0, 3)), 0, 10) -- 4979
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(18,19),( 2, 5)), 0, 10) -- 4980
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(20,21),( 4, 7)), 0, 10) -- 4981
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(22,23),( 6, 9)), 0, 10) -- 4982
,( 3, E,0,0,((20,23),(18,19),( 0, 1),(99,99),(22,23),(12,15)), 0, 10) -- 4983
,( 3, E,0,0,((22,25),(20,21),( 2, 3),(99,99),(24,25),(14,17)), 0, 10) -- 4984
,( 3, E,0,0,((24,27),(22,23),( 4, 5),(99,99),(26,27),(16,19)), 0, 10) -- 4985
,( 3, E,0,0,((26,29),(24,25),( 6, 7),(99,99),(28,29),(18,21)), 0, 10) -- 4986
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(20,21),( 2, 5)), 0, 10) -- 4987
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(22,23),( 4, 7)), 0, 10) -- 4988
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(24,25),( 6, 9)), 0, 10) -- 4989
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(26,27),( 8,11)), 0, 10) -- 4990
,( 3, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(18,19),( 0, 3)), 0,  9) -- 4991
,( 3, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(20,21),( 2, 5)), 0,  9) -- 4992
,( 3, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(22,23),( 4, 7)), 0,  9) -- 4993
,( 3, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(24,25),( 6, 9)), 0,  9) -- 4994
,( 3, E,0,0,((22,23),(20,20),( 0, 0),(17,17),(18,18),( 2, 5)), 0,  9) -- 4995
,( 3, E,0,0,((24,25),(22,22),( 2, 2),(19,19),(20,20),( 4, 7)), 0,  9) -- 4996
,( 3, E,0,0,((26,27),(24,24),( 4, 4),(21,21),(22,22),( 6, 9)), 0,  9) -- 4997
,( 3, E,0,0,((28,29),(26,26),( 6, 6),(23,23),(24,24),( 8,11)), 0,  9) -- 4998
,( 3, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(99,99),( 4, 7)), 0,  9) -- 4999
,( 3, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(99,99),( 6, 9)), 0,  9) -- 5000
,( 3, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(99,99),( 8,11)), 0,  9) -- 5001
,( 3, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(99,99),(10,13)), 0,  9) -- 5002
,( 3, E,0,0,((18,21),(18,19),( 0, 1),(20,21),(99,99),( 6, 9)), 0,  9) -- 5003
,( 3, E,0,0,((20,23),(20,21),( 2, 3),(22,23),(99,99),( 8,11)), 0,  9) -- 5004
,( 3, E,0,0,((22,25),(22,23),( 4, 5),(24,25),(99,99),(10,13)), 0,  9) -- 5005
,( 3, E,0,0,((24,27),(24,25),( 6, 7),(26,27),(99,99),(12,15)), 0,  9) -- 5006
,( 3, E,0,0,((18,21),(18,19),( 0, 1),(99,99),(22,23),( 8,11)), 0,  9) -- 5007
,( 3, E,0,0,((20,23),(20,21),( 2, 3),(99,99),(24,25),(10,13)), 0,  9) -- 5008
,( 3, E,0,0,((22,25),(22,23),( 4, 5),(99,99),(26,27),(12,15)), 0,  9) -- 5009
,( 3, E,0,0,((24,27),(24,25),( 6, 7),(99,99),(28,29),(14,17)), 0,  9) -- 5010
,( 3, E,0,0,((20,23),(20,20),( 1, 1),(20,20),(99,99),(10,13)), 0,  9) -- 5011
,( 3, E,0,0,((22,25),(22,22),( 3, 3),(22,22),(99,99),(12,15)), 0,  9) -- 5012
,( 3, E,0,0,((24,27),(24,24),( 5, 5),(24,24),(99,99),(14,17)), 0,  9) -- 5013
,( 3, E,0,0,((26,29),(26,26),( 7, 7),(26,26),(99,99),(16,19)), 0,  9) -- 5014
,( 3, E,0,0,((22,25),(20,21),( 0, 1),(99,99),(22,23),( 4, 7)), 0,  9) -- 5015
,( 3, E,0,0,((24,27),(22,23),( 2, 3),(99,99),(24,25),( 6, 9)), 0,  9) -- 5016
,( 3, E,0,0,((26,29),(24,25),( 4, 5),(99,99),(26,27),( 8,11)), 0,  9) -- 5017
,( 3, E,0,0,((28,31),(26,27),( 6, 7),(99,99),(28,29),(10,13)), 0,  9) -- 5018
,( 3, E,0,0,((18,21),(18,19),( 0, 1),(99,99),(20,21),( 2, 5)), 0,  9) -- 5019
,( 3, E,0,0,((20,23),(20,21),( 2, 3),(99,99),(22,23),( 4, 7)), 0,  9) -- 5020
,( 3, E,0,0,((22,25),(22,23),( 4, 5),(99,99),(24,25),( 6, 9)), 0,  9) -- 5021
,( 3, E,0,0,((24,27),(24,25),( 6, 7),(99,99),(26,27),( 8,11)), 0,  9) -- 5022
,( 3, E,0,0,((20,23),(20,21),( 1, 1),(99,99),(24,24),(12,15)), 0,  9) -- 5023
,( 3, E,0,0,((22,25),(22,23),( 3, 3),(99,99),(26,26),(14,17)), 0,  9) -- 5024
,( 3, E,0,0,((24,27),(24,25),( 5, 5),(99,99),(28,28),(16,19)), 0,  9) -- 5025
,( 3, E,0,0,((26,29),(26,27),( 7, 7),(99,99),(30,30),(18,21)), 0,  9) -- 5026
,( 3, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(18,19),(99,99)), 0,  9) -- 5027
,( 3, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(20,21),(99,99)), 0,  9) -- 5028
,( 3, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(22,23),(99,99)), 0,  9) -- 5029
,( 3, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(24,25),(99,99)), 0,  9) -- 5030
,( 3, E,0,0,((20,23),(19,19),( 0, 0),(18,19),(99,99),( 8, 9)), 0,  9) -- 5031
,( 3, E,0,0,((22,25),(21,21),( 2, 2),(20,21),(99,99),(10,11)), 0,  9) -- 5032
,( 3, E,0,0,((24,27),(23,23),( 4, 4),(22,23),(99,99),(12,13)), 0,  9) -- 5033
,( 3, E,0,0,((26,29),(25,25),( 6, 6),(24,25),(99,99),(14,15)), 0,  9) -- 5034
,( 3, E,0,0,((24,27),(22,23),( 1, 1),(99,99),(24,24),(13,13)), 0,  9) -- 5035
,( 3, E,0,0,((26,29),(24,25),( 3, 3),(99,99),(26,26),(15,15)), 0,  9) -- 5036
,( 3, E,0,0,((28,31),(26,27),( 5, 5),(99,99),(28,28),(17,17)), 0,  9) -- 5037
,( 3, E,0,0,((30,33),(28,29),( 7, 7),(99,99),(30,30),(19,19)), 0,  9) -- 5038
,( 3, E,0,0,((16,19),(16,17),( 0, 0),(18,19),(99,99),(15,15)), 0,  9) -- 5039
,( 3, E,0,0,((18,21),(18,19),( 2, 2),(20,21),(99,99),(17,17)), 0,  9) -- 5040
,( 3, E,0,0,((20,23),(20,21),( 4, 4),(22,23),(99,99),(19,19)), 0,  9) -- 5041
,( 3, E,0,0,((22,25),(22,23),( 6, 6),(24,25),(99,99),(21,21)), 0,  9) -- 5042
,( 3, E,0,0,((20,23),(19,19),( 0, 0),(99,99),(18,19),( 2, 5)), 0,  9) -- 5043
,( 3, E,0,0,((22,25),(21,21),( 2, 2),(99,99),(20,21),( 4, 7)), 0,  9) -- 5044
,( 3, E,0,0,((24,27),(23,23),( 4, 4),(99,99),(22,23),( 6, 9)), 0,  9) -- 5045
,( 3, E,0,0,((26,29),(25,25),( 6, 6),(99,99),(24,25),( 8,11)), 0,  9) -- 5046
,( 3, E,0,0,((20,23),(19,19),( 0, 1),(18,19),(99,99),( 2, 5)), 0,  9) -- 5047
,( 3, E,0,0,((22,25),(21,21),( 2, 3),(20,21),(99,99),( 4, 7)), 0,  9) -- 5048
,( 3, E,0,0,((24,27),(23,23),( 4, 5),(22,23),(99,99),( 6, 9)), 0,  9) -- 5049
,( 3, E,0,0,((26,29),(25,25),( 6, 7),(24,25),(99,99),( 8,11)), 0,  9) -- 5050
,( 3, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(99,99),( 6, 9)), 0,  9) -- 5051
,( 3, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(99,99),( 8,11)), 0,  9) -- 5052
,( 3, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(99,99),(10,13)), 0,  9) -- 5053
,( 3, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(99,99),(12,15)), 0,  9) -- 5054
,( 3, E,0,0,((20,23),(19,19),( 0, 0),(18,18),(17,17),(99,99)), 0,  9) -- 5055
,( 3, E,0,0,((22,25),(21,21),( 2, 2),(20,20),(19,19),(99,99)), 0,  9) -- 5056
,( 3, E,0,0,((24,27),(23,23),( 4, 4),(22,22),(21,21),(99,99)), 0,  9) -- 5057
,( 3, E,0,0,((26,29),(25,25),( 6, 6),(24,24),(23,23),(99,99)), 0,  9) -- 5058
,( 3, E,0,0,((20,23),(18,19),( 0, 1),(99,99),(21,21),( 4, 7)), 0,  9) -- 5059
,( 3, E,0,0,((22,25),(20,21),( 2, 3),(99,99),(23,23),( 6, 9)), 0,  9) -- 5060
,( 3, E,0,0,((24,27),(22,23),( 4, 5),(99,99),(25,25),( 8,11)), 0,  9) -- 5061
,( 3, E,0,0,((26,29),(24,25),( 6, 7),(99,99),(27,27),(10,13)), 0,  9) -- 5062
,( 3, E,0,0,((21,21),(20,20),( 1, 1),(19,19),(99,99),( 6, 9)), 0,  9) -- 5063
,( 3, E,0,0,((23,23),(22,22),( 3, 3),(21,21),(99,99),( 8,11)), 0,  9) -- 5064
,( 3, E,0,0,((25,25),(24,24),( 5, 5),(23,23),(99,99),(10,13)), 0,  9) -- 5065
,( 3, E,0,0,((27,27),(26,26),( 7, 7),(25,25),(99,99),(12,15)), 0,  9) -- 5066
,( 3, E,0,0,((20,21),(20,20),( 1, 1),(99,99),(22,23),( 4, 7)), 0,  9) -- 5067
,( 3, E,0,0,((22,23),(22,22),( 3, 3),(99,99),(24,25),( 6, 9)), 0,  9) -- 5068
,( 3, E,0,0,((24,25),(24,24),( 5, 5),(99,99),(26,27),( 8,11)), 0,  9) -- 5069
,( 3, E,0,0,((26,27),(26,26),( 7, 7),(99,99),(28,29),(10,13)), 0,  9) -- 5070
,( 3, E,0,0,((25,25),(22,22),( 1, 1),(99,99),(22,23),( 6, 7)), 0,  9) -- 5071
,( 3, E,0,0,((27,27),(24,24),( 3, 3),(99,99),(24,25),( 8, 9)), 0,  9) -- 5072
,( 3, E,0,0,((29,29),(26,26),( 5, 5),(99,99),(26,27),(10,11)), 0,  9) -- 5073
,( 3, E,0,0,((31,31),(28,28),( 7, 7),(99,99),(28,29),(12,13)), 0,  9) -- 5074
,( 3, E,0,0,((18,21),(18,19),( 0, 0),(99,99),(22,22),( 6, 7)), 0,  9) -- 5075
,( 3, E,0,0,((20,23),(20,21),( 2, 2),(99,99),(24,24),( 8, 9)), 0,  9) -- 5076
,( 3, E,0,0,((22,25),(22,23),( 4, 4),(99,99),(26,26),(10,11)), 0,  9) -- 5077
,( 3, E,0,0,((24,27),(24,25),( 6, 6),(99,99),(28,28),(12,13)), 0,  9) -- 5078
,( 3, E,0,0,((18,21),(17,17),( 0, 0),(99,99),(20,21),( 6, 9)), 0,  9) -- 5079
,( 3, E,0,0,((20,23),(19,19),( 2, 2),(99,99),(22,23),( 8,11)), 0,  9) -- 5080
,( 3, E,0,0,((22,25),(21,21),( 4, 4),(99,99),(24,25),(10,13)), 0,  9) -- 5081
,( 3, E,0,0,((24,27),(23,23),( 6, 6),(99,99),(26,27),(12,15)), 0,  9) -- 5082
,( 3, E,0,0,((14,17),(16,19),( 0, 1),(18,21),(18,21),(99,99)), 0,  8) -- 5083
,( 3, E,0,0,((16,19),(18,21),( 2, 3),(20,23),(20,23),(99,99)), 0,  8) -- 5084
,( 3, E,0,0,((18,21),(20,23),( 4, 5),(22,25),(22,25),(99,99)), 0,  8) -- 5085
,( 3, E,0,0,((20,23),(22,25),( 6, 7),(24,27),(24,27),(99,99)), 0,  8) -- 5086
,( 3, E,0,0,((18,21),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 5087
,( 3, E,0,0,((20,23),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 5088
,( 3, E,0,0,((22,25),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 5089
,( 3, E,0,0,((24,27),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 5090
,( 3, E,0,0,((18,21),(18,21),( 0, 1),(18,21),(18,21),(99,99)), 0,  8) -- 5091
,( 3, E,0,0,((20,23),(20,23),( 2, 3),(20,23),(20,23),(99,99)), 0,  8) -- 5092
,( 3, E,0,0,((22,25),(22,25),( 4, 5),(22,25),(22,25),(99,99)), 0,  8) -- 5093
,( 3, E,0,0,((24,27),(24,27),( 6, 7),(24,27),(24,27),(99,99)), 0,  8) -- 5094
,( 3, E,0,0,((22,25),(20,23),( 0, 1),(16,19),(14,17),(99,99)), 0,  7) -- 5095
,( 3, E,0,0,((24,27),(22,25),( 2, 3),(18,21),(16,19),(99,99)), 0,  7) -- 5096
,( 3, E,0,0,((26,29),(24,27),( 4, 5),(20,23),(18,21),(99,99)), 0,  7) -- 5097
,( 3, E,0,0,((28,31),(26,29),( 6, 7),(22,25),(20,23),(99,99)), 0,  7) -- 5098
,( 3, E,0,1,((16,19),(16,19),( 0, 1),(17,17),(99,99),(99,99)), 0,  7) -- 5099
,( 3, E,0,1,((18,21),(18,21),( 2, 3),(19,19),(99,99),(99,99)), 0,  7) -- 5100
,( 3, E,0,1,((20,23),(20,23),( 4, 5),(21,21),(99,99),(99,99)), 0,  7) -- 5101
,( 3, E,0,1,((22,25),(22,25),( 6, 7),(23,23),(99,99),(99,99)), 0,  7) -- 5102
,( 3, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 5103
,( 3, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 5104
,( 3, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 5105
,( 3, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 5106
,( 3, E,0,1,(( 8,11),(12,15),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 5107
,( 3, E,0,1,((10,13),(14,17),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 5108
,( 3, E,0,1,((12,15),(16,19),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 5109
,( 3, E,0,1,((14,17),(18,21),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 5110
,( 3, E,0,1,((12,15),(16,19),( 0, 1),(17,17),(99,99),(99,99)), 0,  6) -- 5111
,( 3, E,0,1,((14,17),(18,21),( 2, 3),(19,19),(99,99),(99,99)), 0,  6) -- 5112
,( 3, E,0,1,((16,19),(20,23),( 4, 5),(21,21),(99,99),(99,99)), 0,  6) -- 5113
,( 3, E,0,1,((18,21),(22,25),( 6, 7),(23,23),(99,99),(99,99)), 0,  6) -- 5114
,( 3, E,0,1,(( 0, 3),(12,13),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 5115
,( 3, E,0,1,(( 2, 5),(14,15),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 5116
,( 3, E,0,1,(( 4, 7),(16,17),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 5117
,( 3, E,0,1,(( 6, 9),(18,19),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 5118
,( 3, E,0,1,((18,21),(20,23),( 0, 1),(99,99),(99,99),(99,99)), 0,  6) -- 5119
,( 3, E,0,1,((20,23),(22,25),( 2, 3),(99,99),(99,99),(99,99)), 0,  6) -- 5120
,( 3, E,0,1,((22,25),(24,27),( 4, 5),(99,99),(99,99),(99,99)), 0,  6) -- 5121
,( 3, E,0,1,((24,27),(26,29),( 6, 7),(99,99),(99,99),(99,99)), 0,  6) -- 5122
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 5123
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 5124
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 5125
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 5126
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 5127
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 5128
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 5129
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 5130
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 5131
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 5132
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 5133
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 5134
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 5135
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 5136
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 5137
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 5138
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(99,99),( 9, 9)), 1, 31) -- 5139
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(99,99),(10,10)), 1, 31) -- 5140
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(99,99),(11,11)), 1, 31) -- 5141
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(99,99),(12,12)), 1, 31) -- 5142
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(99,99),(13,13)), 1, 31) -- 5143
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(99,99),(14,14)), 1, 31) -- 5144
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(99,99),(15,15)), 1, 31) -- 5145
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(99,99),(16,16)), 1, 31) -- 5146
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 30) -- 5147
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 30) -- 5148
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 30) -- 5149
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 30) -- 5150
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 30) -- 5151
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 30) -- 5152
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 30) -- 5153
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 30) -- 5154
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 29) -- 5155
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 29) -- 5156
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 29) -- 5157
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 29) -- 5158
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 29) -- 5159
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 29) -- 5160
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 29) -- 5161
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 29) -- 5162
,( 4, E,0,0,((32,32),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 29) -- 5163
,( 4, E,0,0,((33,33),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 29) -- 5164
,( 4, E,0,0,((34,34),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 1, 29) -- 5165
,( 4, E,0,0,((35,35),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 1, 29) -- 5166
,( 4, E,0,0,((36,36),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 1, 29) -- 5167
,( 4, E,0,0,((37,37),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 1, 29) -- 5168
,( 4, E,0,0,((38,38),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 1, 29) -- 5169
,( 4, E,0,0,((39,39),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 1, 29) -- 5170
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 28) -- 5171
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 28) -- 5172
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 28) -- 5173
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 28) -- 5174
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 28) -- 5175
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 28) -- 5176
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 28) -- 5177
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 28) -- 5178
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 28) -- 5179
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 28) -- 5180
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 28) -- 5181
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 28) -- 5182
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 28) -- 5183
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 28) -- 5184
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 28) -- 5185
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 28) -- 5186
,( 4, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 26) -- 5187
,( 4, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 26) -- 5188
,( 4, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 26) -- 5189
,( 4, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 26) -- 5190
,( 4, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 26) -- 5191
,( 4, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 26) -- 5192
,( 4, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 26) -- 5193
,( 4, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 26) -- 5194
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 25) -- 5195
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 25) -- 5196
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 25) -- 5197
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 25) -- 5198
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 25) -- 5199
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 25) -- 5200
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 25) -- 5201
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 25) -- 5202
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 5203
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 5204
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 5205
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 5206
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 5207
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 5208
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 5209
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 5210
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 5211
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 5212
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 5213
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 5214
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 5215
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 5216
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 5217
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 5218
,( 4, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 23) -- 5219
,( 4, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 23) -- 5220
,( 4, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 23) -- 5221
,( 4, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 23) -- 5222
,( 4, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 23) -- 5223
,( 4, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 23) -- 5224
,( 4, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 23) -- 5225
,( 4, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 23) -- 5226
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 22) -- 5227
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 22) -- 5228
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 22) -- 5229
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 22) -- 5230
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 22) -- 5231
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 22) -- 5232
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 22) -- 5233
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 22) -- 5234
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 21) -- 5235
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 21) -- 5236
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 21) -- 5237
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 21) -- 5238
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 21) -- 5239
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 21) -- 5240
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 21) -- 5241
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 21) -- 5242
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 5243
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 5244
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 5245
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 5246
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 5247
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 5248
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 5249
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 5250
,( 4, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 5251
,( 4, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 5252
,( 4, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 5253
,( 4, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 5254
,( 4, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 5255
,( 4, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 5256
,( 4, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 5257
,( 4, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 5258
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 5259
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 5260
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 5261
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 5262
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 5263
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 5264
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 5265
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 5266
,( 4, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 5267
,( 4, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 5268
,( 4, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 5269
,( 4, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 5270
,( 4, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 5271
,( 4, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 5272
,( 4, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 5273
,( 4, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 5274
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 18) -- 5275
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 18) -- 5276
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 18) -- 5277
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 18) -- 5278
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 18) -- 5279
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 18) -- 5280
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 18) -- 5281
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 18) -- 5282
,( 4, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 5283
,( 4, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 5284
,( 4, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 5285
,( 4, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 5286
,( 4, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 5287
,( 4, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 5288
,( 4, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 5289
,( 4, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 5290
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 5291
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 5292
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 5293
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 5294
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 5295
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 5296
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 5297
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 5298
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 5299
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 5300
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 5301
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 5302
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 5303
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 5304
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 5305
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 5306
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 5307
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 5308
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 5309
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 5310
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 5311
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 5312
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 5313
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 5314
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 5315
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 5316
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 5317
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 5318
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 5319
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 5320
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 5321
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 5322
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 5323
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 5324
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 5325
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 5326
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 5327
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 5328
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 5329
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 5330
,( 4, E,0,0,((34,34),(24,24),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 5331
,( 4, E,0,0,((35,35),(25,25),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 5332
,( 4, E,0,0,((36,36),(26,26),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 5333
,( 4, E,0,0,((37,37),(27,27),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 5334
,( 4, E,0,0,((38,38),(28,28),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 5335
,( 4, E,0,0,((39,39),(29,29),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 5336
,( 4, E,0,0,((40,40),(30,30),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 5337
,( 4, E,0,0,((41,41),(31,31),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 5338
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 5339
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 5340
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 5341
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 5342
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 5343
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 5344
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 5345
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 5346
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 5347
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 5348
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 5349
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 5350
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 5351
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 5352
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 5353
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 5354
,( 4, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 16) -- 5355
,( 4, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 16) -- 5356
,( 4, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 16) -- 5357
,( 4, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 16) -- 5358
,( 4, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 16) -- 5359
,( 4, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 16) -- 5360
,( 4, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 16) -- 5361
,( 4, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 16) -- 5362
,( 4, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 16) -- 5363
,( 4, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 16) -- 5364
,( 4, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 16) -- 5365
,( 4, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 16) -- 5366
,( 4, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 16) -- 5367
,( 4, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 16) -- 5368
,( 4, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 16) -- 5369
,( 4, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 16) -- 5370
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 16) -- 5371
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 16) -- 5372
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 16) -- 5373
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 16) -- 5374
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 16) -- 5375
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 16) -- 5376
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 16) -- 5377
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 16) -- 5378
,( 4, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 5379
,( 4, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 5380
,( 4, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 5381
,( 4, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 5382
,( 4, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 5383
,( 4, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 5384
,( 4, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 5385
,( 4, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 5386
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 5387
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 5388
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 5389
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 5390
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 5391
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 5392
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 5393
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 5394
,( 4, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 5395
,( 4, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 5396
,( 4, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 5397
,( 4, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 5398
,( 4, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 5399
,( 4, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 5400
,( 4, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 5401
,( 4, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 5402
,( 4, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 5403
,( 4, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 5404
,( 4, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 5405
,( 4, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 5406
,( 4, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 5407
,( 4, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 5408
,( 4, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 5409
,( 4, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 5410
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 5411
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 5412
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 5413
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 5414
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 5415
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 5416
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 5417
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 5418
,( 4, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 5419
,( 4, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 5420
,( 4, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 5421
,( 4, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 5422
,( 4, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 5423
,( 4, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 5424
,( 4, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 5425
,( 4, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 5426
,( 4, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 15) -- 5427
,( 4, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 15) -- 5428
,( 4, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 15) -- 5429
,( 4, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 15) -- 5430
,( 4, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 15) -- 5431
,( 4, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 15) -- 5432
,( 4, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 15) -- 5433
,( 4, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 15) -- 5434
,( 4, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 5435
,( 4, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 5436
,( 4, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 5437
,( 4, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 5438
,( 4, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 5439
,( 4, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 5440
,( 4, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 5441
,( 4, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 5442
,( 4, E,0,0,((34,37),(25,25),( 0, 0),(14,15),(14,15),( 4, 7)), 1, 14) -- 5443
,( 4, E,0,0,((36,39),(27,27),( 2, 2),(16,17),(16,17),( 6, 9)), 1, 14) -- 5444
,( 4, E,0,0,((38,41),(29,29),( 4, 4),(18,19),(18,19),( 8,11)), 1, 14) -- 5445
,( 4, E,0,0,((40,43),(31,31),( 6, 6),(20,21),(20,21),(10,13)), 1, 14) -- 5446
,( 4, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 13) -- 5447
,( 4, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),( 8,11)), 1, 13) -- 5448
,( 4, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),(10,13)), 1, 13) -- 5449
,( 4, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(12,15)), 1, 13) -- 5450
,( 4, E,0,0,((36,39),(26,27),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 13) -- 5451
,( 4, E,0,0,((38,41),(28,29),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 13) -- 5452
,( 4, E,0,0,((40,43),(30,31),( 5, 5),(20,20),(18,19),( 8,11)), 1, 13) -- 5453
,( 4, E,0,0,((42,45),(32,33),( 7, 7),(22,22),(20,21),(10,13)), 1, 13) -- 5454
,( 4, E,0,0,((34,37),(25,25),( 0, 0),(14,14),(12,13),( 2, 5)), 1, 13) -- 5455
,( 4, E,0,0,((36,39),(27,27),( 2, 2),(16,16),(14,15),( 4, 7)), 1, 13) -- 5456
,( 4, E,0,0,((38,41),(29,29),( 4, 4),(18,18),(16,17),( 6, 9)), 1, 13) -- 5457
,( 4, E,0,0,((40,43),(31,31),( 6, 6),(20,20),(18,19),( 8,11)), 1, 13) -- 5458
,( 4, E,0,0,((38,41),(28,28),( 1, 1),(15,15),(14,15),( 4, 7)), 1, 12) -- 5459
,( 4, E,0,0,((40,43),(30,30),( 3, 3),(17,17),(16,17),( 6, 9)), 1, 12) -- 5460
,( 4, E,0,0,((42,45),(32,32),( 5, 5),(19,19),(18,19),( 8,11)), 1, 12) -- 5461
,( 4, E,0,0,((44,47),(34,34),( 7, 7),(21,21),(20,21),(10,13)), 1, 12) -- 5462
,( 4, E,0,0,((38,41),(28,28),( 1, 1),(14,15),(13,13),( 4, 7)), 1, 12) -- 5463
,( 4, E,0,0,((40,43),(30,30),( 3, 3),(16,17),(15,15),( 6, 9)), 1, 12) -- 5464
,( 4, E,0,0,((42,45),(32,32),( 5, 5),(18,19),(17,17),( 8,11)), 1, 12) -- 5465
,( 4, E,0,0,((44,47),(34,34),( 7, 7),(20,21),(19,19),(10,13)), 1, 12) -- 5466
,( 4, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 6, 7)), 1, 12) -- 5467
,( 4, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 8, 9)), 1, 12) -- 5468
,( 4, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),(10,11)), 1, 12) -- 5469
,( 4, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),(12,13)), 1, 12) -- 5470
,( 4, E,0,0,((38,38),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 12) -- 5471
,( 4, E,0,0,((40,40),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 12) -- 5472
,( 4, E,0,0,((42,42),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 12) -- 5473
,( 4, E,0,0,((44,44),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 12) -- 5474
,( 4, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 5475
,( 4, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 5476
,( 4, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 5477
,( 4, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 5478
,( 4, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(10,11),( 2, 5)), 1, 11) -- 5479
,( 4, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(12,13),( 4, 7)), 1, 11) -- 5480
,( 4, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(14,15),( 6, 9)), 1, 11) -- 5481
,( 4, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(16,17),( 8,11)), 1, 11) -- 5482
,( 4, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(12,13),( 4, 7)), 1, 11) -- 5483
,( 4, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(14,15),( 6, 9)), 1, 11) -- 5484
,( 4, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(16,17),( 8,11)), 1, 11) -- 5485
,( 4, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(18,19),(10,13)), 1, 11) -- 5486
,( 4, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 8,11)), 1, 11) -- 5487
,( 4, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(10,13)), 1, 11) -- 5488
,( 4, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(12,15)), 1, 11) -- 5489
,( 4, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(14,17)), 1, 11) -- 5490
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 5491
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 5492
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 10) -- 5493
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 10) -- 5494
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 5495
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 5496
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 5497
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 5498
,( 4, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 8,11)), 1, 10) -- 5499
,( 4, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),(10,13)), 1, 10) -- 5500
,( 4, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),(12,15)), 1, 10) -- 5501
,( 4, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),(14,17)), 1, 10) -- 5502
,( 4, E,0,0,((38,41),(26,27),( 0, 1),(14,15),(14,15),(10,13)), 1, 10) -- 5503
,( 4, E,0,0,((40,43),(28,29),( 2, 3),(16,17),(16,17),(12,15)), 1, 10) -- 5504
,( 4, E,0,0,((42,45),(30,31),( 4, 5),(18,19),(18,19),(14,17)), 1, 10) -- 5505
,( 4, E,0,0,((44,47),(32,33),( 6, 7),(20,21),(20,21),(16,19)), 1, 10) -- 5506
,( 4, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),(12,15)), 1, 10) -- 5507
,( 4, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(14,17)), 1, 10) -- 5508
,( 4, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(16,19)), 1, 10) -- 5509
,( 4, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(18,21)), 1, 10) -- 5510
,( 4, E,0,0,((40,40),(27,27),( 0, 0),(13,13),(10,11),( 2, 5)), 1, 10) -- 5511
,( 4, E,0,0,((42,42),(29,29),( 2, 2),(15,15),(12,13),( 4, 7)), 1, 10) -- 5512
,( 4, E,0,0,((44,44),(31,31),( 4, 4),(17,17),(14,15),( 6, 9)), 1, 10) -- 5513
,( 4, E,0,0,((46,46),(33,33),( 6, 6),(19,19),(16,17),( 8,11)), 1, 10) -- 5514
,( 4, E,0,0,((38,41),(26,27),( 0, 0),(13,13),(12,13),( 6, 9)), 1, 10) -- 5515
,( 4, E,0,0,((40,43),(28,29),( 2, 2),(15,15),(14,15),( 8,11)), 1, 10) -- 5516
,( 4, E,0,0,((42,45),(30,31),( 4, 4),(17,17),(16,17),(10,13)), 1, 10) -- 5517
,( 4, E,0,0,((44,47),(32,33),( 6, 6),(19,19),(18,19),(12,15)), 1, 10) -- 5518
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(10,11),( 0, 1)), 1, 10) -- 5519
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(12,13),( 2, 3)), 1, 10) -- 5520
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(14,15),( 4, 5)), 1, 10) -- 5521
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(16,17),( 6, 7)), 1, 10) -- 5522
,( 4, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(15,15),(14,15)), 1, 10) -- 5523
,( 4, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(17,17),(16,17)), 1, 10) -- 5524
,( 4, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(19,19),(18,19)), 1, 10) -- 5525
,( 4, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(21,21),(20,21)), 1, 10) -- 5526
,( 4, E,0,0,((38,41),(28,28),( 0, 1),(99,99),(13,13),( 8,11)), 1, 10) -- 5527
,( 4, E,0,0,((40,43),(30,30),( 2, 3),(99,99),(15,15),(10,13)), 1, 10) -- 5528
,( 4, E,0,0,((42,45),(32,32),( 4, 5),(99,99),(17,17),(12,15)), 1, 10) -- 5529
,( 4, E,0,0,((44,47),(34,34),( 6, 7),(99,99),(19,19),(14,17)), 1, 10) -- 5530
,( 4, E,0,0,((40,41),(28,29),( 0, 1),(99,99),( 8, 9),( 0, 1)), 1, 10) -- 5531
,( 4, E,0,0,((42,43),(30,31),( 2, 3),(99,99),(10,11),( 2, 3)), 1, 10) -- 5532
,( 4, E,0,0,((44,45),(32,33),( 4, 5),(99,99),(12,13),( 4, 5)), 1, 10) -- 5533
,( 4, E,0,0,((46,47),(34,35),( 6, 7),(99,99),(14,15),( 6, 7)), 1, 10) -- 5534
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(14,15),(14,17)), 1,  9) -- 5535
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(16,17),(16,19)), 1,  9) -- 5536
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(18,19),(18,21)), 1,  9) -- 5537
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(20,21),(20,23)), 1,  9) -- 5538
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(15,15),(16,17),(14,17)), 1,  9) -- 5539
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(17,17),(18,19),(16,19)), 1,  9) -- 5540
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(19,19),(20,21),(18,21)), 1,  9) -- 5541
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(21,21),(22,23),(20,23)), 1,  9) -- 5542
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(10,11),( 6, 9)), 1,  9) -- 5543
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(12,13),( 8,11)), 1,  9) -- 5544
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(14,15),(10,13)), 1,  9) -- 5545
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(16,17),(12,15)), 1,  9) -- 5546
,( 4, E,0,0,((38,41),(26,27),( 0, 1),(14,14),(12,13),(10,13)), 1,  9) -- 5547
,( 4, E,0,0,((40,43),(28,29),( 2, 3),(16,16),(14,15),(12,15)), 1,  9) -- 5548
,( 4, E,0,0,((42,45),(30,31),( 4, 5),(18,18),(16,17),(14,17)), 1,  9) -- 5549
,( 4, E,0,0,((44,47),(32,33),( 6, 7),(20,20),(18,19),(16,19)), 1,  9) -- 5550
,( 4, E,0,0,((42,42),(29,29),( 1, 1),(15,15),(14,14),( 8,11)), 1,  9) -- 5551
,( 4, E,0,0,((44,44),(31,31),( 3, 3),(17,17),(16,16),(10,13)), 1,  9) -- 5552
,( 4, E,0,0,((46,46),(33,33),( 5, 5),(19,19),(18,18),(12,15)), 1,  9) -- 5553
,( 4, E,0,0,((48,48),(35,35),( 7, 7),(21,21),(20,20),(14,17)), 1,  9) -- 5554
,( 4, E,0,0,((40,40),(27,27),( 0, 0),(13,13),(11,11),( 6, 9)), 1,  9) -- 5555
,( 4, E,0,0,((42,42),(29,29),( 2, 2),(15,15),(13,13),( 8,11)), 1,  9) -- 5556
,( 4, E,0,0,((44,44),(31,31),( 4, 4),(17,17),(15,15),(10,13)), 1,  9) -- 5557
,( 4, E,0,0,((46,46),(33,33),( 6, 6),(19,19),(17,17),(12,15)), 1,  9) -- 5558
,( 4, E,0,0,((41,41),(28,28),( 1, 1),(15,15),(14,15),(18,21)), 1,  9) -- 5559
,( 4, E,0,0,((43,43),(30,30),( 3, 3),(17,17),(16,17),(20,23)), 1,  9) -- 5560
,( 4, E,0,0,((45,45),(32,32),( 5, 5),(19,19),(18,19),(22,23)), 1,  9) -- 5561
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(99,99),(12,13),(10,13)), 1,  9) -- 5562
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(99,99),(14,15),(12,15)), 1,  9) -- 5563
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(99,99),(16,17),(14,17)), 1,  9) -- 5564
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(99,99),(18,19),(16,19)), 1,  9) -- 5565
,( 4, E,0,0,((40,41),(28,29),( 0, 1),(99,99),(13,13),(14,17)), 1,  9) -- 5566
,( 4, E,0,0,((42,43),(30,31),( 2, 3),(99,99),(15,15),(16,19)), 1,  9) -- 5567
,( 4, E,0,0,((44,45),(32,33),( 4, 5),(99,99),(17,17),(18,21)), 1,  9) -- 5568
,( 4, E,0,0,((46,47),(34,35),( 6, 7),(99,99),(19,19),(20,23)), 1,  9) -- 5569
,( 4, E,0,0,((40,43),(28,29),( 0, 1),(99,99),( 8, 9),( 4, 7)), 1,  9) -- 5570
,( 4, E,0,0,((42,45),(30,31),( 2, 3),(99,99),(10,11),( 6, 9)), 1,  9) -- 5571
,( 4, E,0,0,((44,47),(32,33),( 4, 5),(99,99),(12,13),( 8,11)), 1,  9) -- 5572
,( 4, E,0,0,((46,49),(34,35),( 6, 7),(99,99),(14,15),(10,13)), 1,  9) -- 5573
,( 4, E,0,0,((43,43),(30,30),( 1, 1),(99,99),(12,13),( 8,11)), 1,  9) -- 5574
,( 4, E,0,0,((45,45),(32,32),( 3, 3),(99,99),(14,15),(10,13)), 1,  9) -- 5575
,( 4, E,0,0,((47,47),(34,34),( 5, 5),(99,99),(16,17),(12,15)), 1,  9) -- 5576
,( 4, E,0,0,((49,49),(36,36),( 7, 7),(99,99),(18,19),(14,17)), 1,  9) -- 5577
,( 4, E,0,0,((43,43),(30,30),( 1, 1),(99,99),(10,11),( 4, 7)), 1,  9) -- 5578
,( 4, E,0,0,((45,45),(32,32),( 3, 3),(99,99),(12,13),( 6, 9)), 1,  9) -- 5579
,( 4, E,0,0,((47,47),(34,34),( 5, 5),(99,99),(14,15),( 8,11)), 1,  9) -- 5580
,( 4, E,0,0,((49,49),(36,36),( 7, 7),(99,99),(16,17),(10,13)), 1,  9) -- 5581
,( 4, E,0,0,((46,49),(99,99),( 0, 1),(12,13),(10,11),( 5, 5)), 1,  9) -- 5582
,( 4, E,0,0,((48,51),(99,99),( 2, 3),(14,15),(12,13),( 7, 7)), 1,  9) -- 5583
,( 4, E,0,0,((50,53),(99,99),( 4, 5),(16,17),(14,15),( 9, 9)), 1,  9) -- 5584
,( 4, E,0,0,((52,55),(99,99),( 6, 7),(18,19),(16,17),(11,11)), 1,  9) -- 5585
,( 4, E,0,0,((42,42),(29,29),( 1, 1),(99,99),(14,14),(12,12)), 1,  9) -- 5586
,( 4, E,0,0,((44,44),(31,31),( 3, 3),(99,99),(16,16),(14,14)), 1,  9) -- 5587
,( 4, E,0,0,((46,46),(33,33),( 5, 5),(99,99),(18,18),(16,16)), 1,  9) -- 5588
,( 4, E,0,0,((48,48),(35,35),( 7, 7),(99,99),(20,20),(18,18)), 1,  9) -- 5589
,( 4, E,0,0,((40,43),(28,29),( 0, 0),(99,99),(11,11),(10,13)), 1,  9) -- 5590
,( 4, E,0,0,((42,45),(30,31),( 2, 2),(99,99),(13,13),(12,15)), 1,  9) -- 5591
,( 4, E,0,0,((44,47),(32,33),( 4, 4),(99,99),(15,15),(14,17)), 1,  9) -- 5592
,( 4, E,0,0,((46,49),(34,35),( 6, 6),(99,99),(17,17),(16,19)), 1,  9) -- 5593
,( 4, E,0,0,((48,48),(99,99),( 0, 1),(12,13),( 8, 9),( 4, 4)), 1,  9) -- 5594
,( 4, E,0,0,((50,50),(99,99),( 2, 3),(14,15),(10,11),( 6, 6)), 1,  9) -- 5595
,( 4, E,0,0,((52,52),(99,99),( 4, 5),(16,17),(12,13),( 8, 8)), 1,  9) -- 5596
,( 4, E,0,0,((54,54),(99,99),( 6, 7),(18,19),(14,15),(10,10)), 1,  9) -- 5597
,( 4, E,0,0,((42,45),(30,30),( 1, 1),(99,99),(14,15),(99,99)), 1,  9) -- 5598
,( 4, E,0,0,((44,47),(32,32),( 3, 3),(99,99),(16,17),(99,99)), 1,  9) -- 5599
,( 4, E,0,0,((46,49),(34,34),( 5, 5),(99,99),(18,19),(99,99)), 1,  9) -- 5600
,( 4, E,0,0,((48,51),(36,36),( 7, 7),(99,99),(20,21),(99,99)), 1,  9) -- 5601
,( 4, E,0,0,((40,43),(28,31),( 1, 1),(14,17),(14,17),(99,99)), 1,  8) -- 5602
,( 4, E,0,0,((42,45),(30,33),( 3, 3),(16,19),(16,19),(99,99)), 1,  8) -- 5603
,( 4, E,0,0,((44,47),(32,35),( 5, 5),(18,21),(18,21),(99,99)), 1,  8) -- 5604
,( 4, E,0,0,((46,49),(34,37),( 7, 7),(20,23),(20,23),(99,99)), 1,  8) -- 5605
,( 4, E,0,0,((46,49),(99,99),( 0, 1),(10,13),( 8,11),(99,99)), 1,  8) -- 5606
,( 4, E,0,0,((48,51),(99,99),( 2, 3),(12,15),(10,13),(99,99)), 1,  8) -- 5607
,( 4, E,0,0,((50,53),(99,99),( 4, 5),(14,17),(12,15),(99,99)), 1,  8) -- 5608
,( 4, E,0,0,((52,55),(99,99),( 6, 7),(16,19),(14,17),(99,99)), 1,  8) -- 5609
,( 4, E,0,0,((50,51),(99,99),( 0, 1),(12,13),(10,13),(99,99)), 1,  8) -- 5610
,( 4, E,0,0,((52,53),(99,99),( 2, 3),(14,15),(12,15),(99,99)), 1,  8) -- 5611
,( 4, E,0,0,((54,55),(99,99),( 4, 5),(16,17),(14,17),(99,99)), 1,  8) -- 5612
,( 4, E,0,0,((56,57),(99,99),( 6, 7),(18,19),(16,19),(99,99)), 1,  8) -- 5613
,( 4, E,0,1,((44,47),(28,31),( 0, 1),(14,17),(99,99),(99,99)), 1,  7) -- 5614
,( 4, E,0,1,((46,49),(30,33),( 2, 3),(16,19),(99,99),(99,99)), 1,  7) -- 5615
,( 4, E,0,1,((48,51),(32,35),( 4, 5),(18,21),(99,99),(99,99)), 1,  7) -- 5616
,( 4, E,0,1,((50,53),(34,37),( 6, 7),(20,23),(99,99),(99,99)), 1,  7) -- 5617
,( 4, E,0,1,((40,43),(26,29),( 0, 1),(14,17),(99,99),(99,99)), 1,  7) -- 5618
,( 4, E,0,1,((42,45),(28,31),( 2, 3),(16,19),(99,99),(99,99)), 1,  7) -- 5619
,( 4, E,0,1,((44,47),(30,33),( 4, 5),(18,21),(99,99),(99,99)), 1,  7) -- 5620
,( 4, E,0,1,((46,49),(32,35),( 6, 7),(20,23),(99,99),(99,99)), 1,  7) -- 5621
,( 4, E,0,1,((48,51),(99,99),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 5622
,( 4, E,0,1,((50,53),(99,99),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 5623
,( 4, E,0,1,((52,55),(99,99),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 5624
,( 4, E,0,1,((54,57),(99,99),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 5625
,( 4, E,0,1,((52,55),(99,99),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 5626
,( 4, E,0,1,((54,57),(99,99),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 5627
,( 4, E,0,1,((56,59),(99,99),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 5628
,( 4, E,0,1,((58,61),(99,99),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 5629
,( 4, E,0,1,((46,49),(99,99),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 5630
,( 4, E,0,1,((48,51),(99,99),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 5631
,( 4, E,0,1,((50,53),(99,99),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 5632
,( 4, E,0,1,((52,55),(99,99),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 5633
,( 4, E,0,1,((48,51),(99,99),( 0, 1),(16,16),(99,99),(99,99)), 1,  7) -- 5634
,( 4, E,0,1,((50,53),(99,99),( 2, 3),(18,18),(99,99),(99,99)), 1,  7) -- 5635
,( 4, E,0,1,((52,55),(99,99),( 4, 5),(20,20),(99,99),(99,99)), 1,  7) -- 5636
,( 4, E,0,1,((54,57),(99,99),( 6, 7),(22,22),(99,99),(99,99)), 1,  7) -- 5637
,( 4, E,0,1,((36,39),(24,27),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 5638
,( 4, E,0,1,((38,41),(26,29),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 5639
,( 4, E,0,1,((40,43),(28,31),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 5640
,( 4, E,0,1,((42,45),(30,33),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 5641
,( 4, E,0,1,((40,43),(26,29),( 1, 1),(18,21),(99,99),(99,99)), 1,  6) -- 5642
,( 4, E,0,1,((42,45),(28,31),( 3, 3),(20,23),(99,99),(99,99)), 1,  6) -- 5643
,( 4, E,0,1,((44,47),(30,33),( 5, 5),(22,25),(99,99),(99,99)), 1,  6) -- 5644
,( 4, E,0,1,((46,49),(32,35),( 7, 7),(24,27),(99,99),(99,99)), 1,  6) -- 5645
,( 4, E,0,1,((50,53),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 5646
,( 4, E,0,1,((52,55),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 5647
,( 4, E,0,1,((54,57),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 5648
,( 4, E,0,1,((56,59),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 5649
,( 4, E,0,1,((46,49),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 5650
,( 4, E,0,1,((48,51),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 5651
,( 4, E,0,1,((50,53),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 5652
,( 4, E,0,1,((52,55),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 5653
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 5654
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 5655
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 5656
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 5657
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 5658
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 5659
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 5660
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 5661
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(99,99),( 8, 8)), 0, 31) -- 5662
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(99,99),( 9, 9)), 0, 31) -- 5663
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(99,99),(10,10)), 0, 31) -- 5664
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(99,99),(11,11)), 0, 31) -- 5665
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(99,99),(12,12)), 0, 31) -- 5666
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(99,99),(13,13)), 0, 31) -- 5667
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(99,99),(14,14)), 0, 31) -- 5668
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(99,99),(15,15)), 0, 31) -- 5669
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 30) -- 5670
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 30) -- 5671
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 30) -- 5672
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 30) -- 5673
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 30) -- 5674
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 30) -- 5675
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 30) -- 5676
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 30) -- 5677
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 29) -- 5678
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 29) -- 5679
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 29) -- 5680
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 29) -- 5681
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 29) -- 5682
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 29) -- 5683
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 29) -- 5684
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 29) -- 5685
,( 4, E,0,0,((32,32),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 29) -- 5686
,( 4, E,0,0,((33,33),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 29) -- 5687
,( 4, E,0,0,((34,34),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 29) -- 5688
,( 4, E,0,0,((35,35),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 29) -- 5689
,( 4, E,0,0,((36,36),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 29) -- 5690
,( 4, E,0,0,((37,37),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 29) -- 5691
,( 4, E,0,0,((38,38),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 29) -- 5692
,( 4, E,0,0,((39,39),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 29) -- 5693
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(99,99),( 8, 8)), 0, 29) -- 5694
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(99,99),( 9, 9)), 0, 29) -- 5695
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(99,99),(10,10)), 0, 29) -- 5696
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(99,99),(11,11)), 0, 29) -- 5697
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(99,99),(12,12)), 0, 29) -- 5698
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(99,99),(13,13)), 0, 29) -- 5699
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(99,99),(14,14)), 0, 29) -- 5700
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(99,99),(15,15)), 0, 29) -- 5701
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 27) -- 5702
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 27) -- 5703
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 27) -- 5704
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 27) -- 5705
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 27) -- 5706
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 27) -- 5707
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 27) -- 5708
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 27) -- 5709
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 26) -- 5710
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 26) -- 5711
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 26) -- 5712
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 26) -- 5713
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 26) -- 5714
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 26) -- 5715
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 26) -- 5716
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 26) -- 5717
,( 4, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 25) -- 5718
,( 4, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 25) -- 5719
,( 4, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 25) -- 5720
,( 4, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 25) -- 5721
,( 4, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 25) -- 5722
,( 4, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 25) -- 5723
,( 4, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 25) -- 5724
,( 4, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 25) -- 5725
,( 4, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 24) -- 5726
,( 4, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 24) -- 5727
,( 4, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 24) -- 5728
,( 4, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 24) -- 5729
,( 4, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 24) -- 5730
,( 4, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 24) -- 5731
,( 4, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 24) -- 5732
,( 4, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 24) -- 5733
,( 4, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 23) -- 5734
,( 4, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 23) -- 5735
,( 4, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 23) -- 5736
,( 4, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 23) -- 5737
,( 4, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 23) -- 5738
,( 4, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 23) -- 5739
,( 4, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 23) -- 5740
,( 4, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 23) -- 5741
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 22) -- 5742
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 22) -- 5743
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 22) -- 5744
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 22) -- 5745
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 22) -- 5746
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 22) -- 5747
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 22) -- 5748
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 22) -- 5749
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 21) -- 5750
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 21) -- 5751
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 21) -- 5752
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 21) -- 5753
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 21) -- 5754
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 21) -- 5755
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 21) -- 5756
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 21) -- 5757
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 20) -- 5758
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 20) -- 5759
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 20) -- 5760
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 20) -- 5761
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 20) -- 5762
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 20) -- 5763
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 20) -- 5764
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 20) -- 5765
,( 4, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 5766
,( 4, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 5767
,( 4, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 5768
,( 4, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 5769
,( 4, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 5770
,( 4, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 5771
,( 4, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 5772
,( 4, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 5773
,( 4, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 5774
,( 4, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 5775
,( 4, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 5776
,( 4, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 5777
,( 4, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 5778
,( 4, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 5779
,( 4, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 5780
,( 4, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 5781
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(17,17),(99,99),(10,10)), 0, 19) -- 5782
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(18,18),(99,99),(11,11)), 0, 19) -- 5783
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(19,19),(99,99),(12,12)), 0, 19) -- 5784
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(20,20),(99,99),(13,13)), 0, 19) -- 5785
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(21,21),(99,99),(14,14)), 0, 19) -- 5786
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(22,22),(99,99),(15,15)), 0, 19) -- 5787
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(23,23),(99,99),(16,16)), 0, 19) -- 5788
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(24,24),(99,99),(17,17)), 0, 19) -- 5789
,( 4, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(99,99),(10,10)), 0, 19) -- 5790
,( 4, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(99,99),(11,11)), 0, 19) -- 5791
,( 4, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(99,99),(12,12)), 0, 19) -- 5792
,( 4, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(99,99),(13,13)), 0, 19) -- 5793
,( 4, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(99,99),(14,14)), 0, 19) -- 5794
,( 4, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(99,99),(15,15)), 0, 19) -- 5795
,( 4, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(99,99),(16,16)), 0, 19) -- 5796
,( 4, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(99,99),(17,17)), 0, 19) -- 5797
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 5798
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 5799
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 5800
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 5801
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 5802
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 5803
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 5804
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 5805
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 18) -- 5806
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 18) -- 5807
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 18) -- 5808
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 18) -- 5809
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 18) -- 5810
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 18) -- 5811
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 18) -- 5812
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 18) -- 5813
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(99,99),(10,10)), 0, 18) -- 5814
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(99,99),(11,11)), 0, 18) -- 5815
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(99,99),(12,12)), 0, 18) -- 5816
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(99,99),(13,13)), 0, 18) -- 5817
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(99,99),(14,14)), 0, 18) -- 5818
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(99,99),(15,15)), 0, 18) -- 5819
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(99,99),(16,16)), 0, 18) -- 5820
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(99,99),(17,17)), 0, 18) -- 5821
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(99,99),(11,11)), 0, 18) -- 5822
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(99,99),(12,12)), 0, 18) -- 5823
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(99,99),(13,13)), 0, 18) -- 5824
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(99,99),(14,14)), 0, 18) -- 5825
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(99,99),(15,15)), 0, 18) -- 5826
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(99,99),(16,16)), 0, 18) -- 5827
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(99,99),(17,17)), 0, 18) -- 5828
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(99,99),(18,18)), 0, 18) -- 5829
,( 4, E,0,0,((31,31),(23,23),( 0, 0),(17,17),(99,99),(11,11)), 0, 18) -- 5830
,( 4, E,0,0,((32,32),(24,24),( 1, 1),(18,18),(99,99),(12,12)), 0, 18) -- 5831
,( 4, E,0,0,((33,33),(25,25),( 2, 2),(19,19),(99,99),(13,13)), 0, 18) -- 5832
,( 4, E,0,0,((34,34),(26,26),( 3, 3),(20,20),(99,99),(14,14)), 0, 18) -- 5833
,( 4, E,0,0,((35,35),(27,27),( 4, 4),(21,21),(99,99),(15,15)), 0, 18) -- 5834
,( 4, E,0,0,((36,36),(28,28),( 5, 5),(22,22),(99,99),(16,16)), 0, 18) -- 5835
,( 4, E,0,0,((37,37),(29,29),( 6, 6),(23,23),(99,99),(17,17)), 0, 18) -- 5836
,( 4, E,0,0,((38,38),(30,30),( 7, 7),(24,24),(99,99),(18,18)), 0, 18) -- 5837
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(99,99),(11,11)), 0, 17) -- 5838
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(99,99),(12,12)), 0, 17) -- 5839
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(99,99),(13,13)), 0, 17) -- 5840
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(99,99),(14,14)), 0, 17) -- 5841
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(99,99),(15,15)), 0, 17) -- 5842
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(99,99),(16,16)), 0, 17) -- 5843
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(99,99),(17,17)), 0, 17) -- 5844
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(99,99),(18,18)), 0, 17) -- 5845
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(99,99),( 9, 9)), 0, 17) -- 5846
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(99,99),(10,10)), 0, 17) -- 5847
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(99,99),(11,11)), 0, 17) -- 5848
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(99,99),(12,12)), 0, 17) -- 5849
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(99,99),(13,13)), 0, 17) -- 5850
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(99,99),(14,14)), 0, 17) -- 5851
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(99,99),(15,15)), 0, 17) -- 5852
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(99,99),(16,16)), 0, 17) -- 5853
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 16) -- 5854
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 16) -- 5855
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 16) -- 5856
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 16) -- 5857
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 16) -- 5858
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 16) -- 5859
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 16) -- 5860
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 16) -- 5861
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 5862
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 5863
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 5864
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 5865
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 5866
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 5867
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 5868
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 5869
,( 4, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 5870
,( 4, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 5871
,( 4, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 5872
,( 4, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 5873
,( 4, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 5874
,( 4, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 5875
,( 4, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 5876
,( 4, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 5877
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(99,99),(11,11)), 0, 16) -- 5878
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(99,99),(12,12)), 0, 16) -- 5879
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(99,99),(13,13)), 0, 16) -- 5880
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(99,99),(14,14)), 0, 16) -- 5881
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(99,99),(15,15)), 0, 16) -- 5882
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(99,99),(16,16)), 0, 16) -- 5883
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(99,99),(17,17)), 0, 16) -- 5884
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(99,99),(18,18)), 0, 16) -- 5885
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(99,99),(10,10)), 0, 16) -- 5886
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(99,99),(11,11)), 0, 16) -- 5887
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(99,99),(12,12)), 0, 16) -- 5888
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(99,99),(13,13)), 0, 16) -- 5889
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(99,99),(14,14)), 0, 16) -- 5890
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(99,99),(15,15)), 0, 16) -- 5891
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(99,99),(16,16)), 0, 16) -- 5892
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(99,99),(17,17)), 0, 16) -- 5893
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(99,99),(10,10)), 0, 16) -- 5894
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(99,99),(11,11)), 0, 16) -- 5895
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(99,99),(12,12)), 0, 16) -- 5896
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(99,99),(13,13)), 0, 16) -- 5897
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(99,99),(14,14)), 0, 16) -- 5898
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(99,99),(15,15)), 0, 16) -- 5899
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(99,99),(16,16)), 0, 16) -- 5900
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(99,99),(17,17)), 0, 16) -- 5901
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(99,99),( 9, 9)), 0, 16) -- 5902
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(99,99),(10,10)), 0, 16) -- 5903
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(99,99),(11,11)), 0, 16) -- 5904
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(99,99),(12,12)), 0, 16) -- 5905
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(99,99),(13,13)), 0, 16) -- 5906
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(99,99),(14,14)), 0, 16) -- 5907
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(99,99),(15,15)), 0, 16) -- 5908
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(99,99),(16,16)), 0, 16) -- 5909
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 5910
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 5911
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 5912
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 5913
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 5914
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 5915
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 5916
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 5917
,( 4, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(99,99),(11,11)), 0, 15) -- 5918
,( 4, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(99,99),(12,12)), 0, 15) -- 5919
,( 4, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(99,99),(13,13)), 0, 15) -- 5920
,( 4, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(99,99),(14,14)), 0, 15) -- 5921
,( 4, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(99,99),(15,15)), 0, 15) -- 5922
,( 4, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(99,99),(16,16)), 0, 15) -- 5923
,( 4, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(99,99),(17,17)), 0, 15) -- 5924
,( 4, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(99,99),(18,18)), 0, 15) -- 5925
,( 4, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(99,99),(10,10)), 0, 15) -- 5926
,( 4, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(99,99),(11,11)), 0, 15) -- 5927
,( 4, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(99,99),(12,12)), 0, 15) -- 5928
,( 4, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(99,99),(13,13)), 0, 15) -- 5929
,( 4, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(99,99),(14,14)), 0, 15) -- 5930
,( 4, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(99,99),(15,15)), 0, 15) -- 5931
,( 4, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(99,99),(16,16)), 0, 15) -- 5932
,( 4, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(99,99),(17,17)), 0, 15) -- 5933
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(99,99),(10,10)), 0, 15) -- 5934
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(99,99),(11,11)), 0, 15) -- 5935
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(99,99),(12,12)), 0, 15) -- 5936
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(99,99),(13,13)), 0, 15) -- 5937
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(99,99),(14,14)), 0, 15) -- 5938
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(99,99),(15,15)), 0, 15) -- 5939
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(99,99),(16,16)), 0, 15) -- 5940
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(99,99),(17,17)), 0, 15) -- 5941
,( 4, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(99,99),(11,11)), 0, 15) -- 5942
,( 4, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(99,99),(12,12)), 0, 15) -- 5943
,( 4, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(99,99),(13,13)), 0, 15) -- 5944
,( 4, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(99,99),(14,14)), 0, 15) -- 5945
,( 4, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(99,99),(15,15)), 0, 15) -- 5946
,( 4, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(99,99),(16,16)), 0, 15) -- 5947
,( 4, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(99,99),(17,17)), 0, 15) -- 5948
,( 4, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(99,99),(18,18)), 0, 15) -- 5949
,( 4, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(99,99),(12,12)), 0, 15) -- 5950
,( 4, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(99,99),(13,13)), 0, 15) -- 5951
,( 4, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(99,99),(14,14)), 0, 15) -- 5952
,( 4, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(99,99),(15,15)), 0, 15) -- 5953
,( 4, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(99,99),(16,16)), 0, 15) -- 5954
,( 4, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(99,99),(17,17)), 0, 15) -- 5955
,( 4, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(99,99),(18,18)), 0, 15) -- 5956
,( 4, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(99,99),(19,19)), 0, 15) -- 5957
,( 4, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(99,99),( 9, 9)), 0, 15) -- 5958
,( 4, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(99,99),(10,10)), 0, 15) -- 5959
,( 4, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(99,99),(11,11)), 0, 15) -- 5960
,( 4, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(99,99),(12,12)), 0, 15) -- 5961
,( 4, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(99,99),(13,13)), 0, 15) -- 5962
,( 4, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(99,99),(14,14)), 0, 15) -- 5963
,( 4, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(99,99),(15,15)), 0, 15) -- 5964
,( 4, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(99,99),(16,16)), 0, 15) -- 5965
,( 4, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(99,99),(11,11)), 0, 15) -- 5966
,( 4, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(99,99),(12,12)), 0, 15) -- 5967
,( 4, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(99,99),(13,13)), 0, 15) -- 5968
,( 4, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(99,99),(14,14)), 0, 15) -- 5969
,( 4, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(99,99),(15,15)), 0, 15) -- 5970
,( 4, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(99,99),(16,16)), 0, 15) -- 5971
,( 4, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(99,99),(17,17)), 0, 15) -- 5972
,( 4, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(99,99),(18,18)), 0, 15) -- 5973
,( 4, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(19,19),(10,13)), 0, 14) -- 5974
,( 4, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(21,21),(12,15)), 0, 14) -- 5975
,( 4, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(23,23),(14,17)), 0, 14) -- 5976
,( 4, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(25,25),(16,19)), 0, 14) -- 5977
,( 4, E,0,0,((28,31),(22,23),( 0, 1),(18,19),(20,21),(12,15)), 0, 14) -- 5978
,( 4, E,0,0,((30,33),(24,25),( 2, 3),(20,21),(22,23),(14,17)), 0, 14) -- 5979
,( 4, E,0,0,((32,35),(26,27),( 4, 5),(22,23),(24,25),(16,19)), 0, 14) -- 5980
,( 4, E,0,0,((34,37),(28,29),( 6, 7),(24,25),(26,27),(18,21)), 0, 14) -- 5981
,( 4, E,0,0,((26,29),(21,21),( 0, 0),(16,17),(20,20),(10,13)), 0, 14) -- 5982
,( 4, E,0,0,((28,31),(23,23),( 2, 2),(18,19),(22,22),(12,15)), 0, 14) -- 5983
,( 4, E,0,0,((30,33),(25,25),( 4, 4),(20,21),(24,24),(14,17)), 0, 14) -- 5984
,( 4, E,0,0,((32,35),(27,27),( 6, 6),(22,23),(26,26),(16,19)), 0, 14) -- 5985
,( 4, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,20),(10,13)), 0, 13) -- 5986
,( 4, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,22),(12,15)), 0, 13) -- 5987
,( 4, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,24),(14,17)), 0, 13) -- 5988
,( 4, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,26),(16,19)), 0, 13) -- 5989
,( 4, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 5990
,( 4, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 5991
,( 4, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 5992
,( 4, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 5993
,( 4, E,0,0,((26,27),(22,22),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 5994
,( 4, E,0,0,((28,29),(24,24),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 5995
,( 4, E,0,0,((30,31),(26,26),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 5996
,( 4, E,0,0,((32,33),(28,28),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 5997
,( 4, E,0,0,((24,27),(20,21),( 0, 0),(16,17),(19,19),( 8,11)), 0, 12) -- 5998
,( 4, E,0,0,((26,29),(22,23),( 2, 2),(18,19),(21,21),(10,13)), 0, 12) -- 5999
,( 4, E,0,0,((28,31),(24,25),( 4, 4),(20,21),(23,23),(12,15)), 0, 12) -- 6000
,( 4, E,0,0,((30,33),(26,27),( 6, 6),(22,23),(25,25),(14,17)), 0, 12) -- 6001
,( 4, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(12,15)), 0, 12) -- 6002
,( 4, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(14,17)), 0, 12) -- 6003
,( 4, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(16,19)), 0, 12) -- 6004
,( 4, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(18,21)), 0, 12) -- 6005
,( 4, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(22,23),(14,17)), 0, 12) -- 6006
,( 4, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(24,25),(16,19)), 0, 12) -- 6007
,( 4, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(26,27),(18,21)), 0, 12) -- 6008
,( 4, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(28,29),(20,23)), 0, 12) -- 6009
,( 4, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(20,20),(10,13)), 0, 12) -- 6010
,( 4, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(22,22),(12,15)), 0, 12) -- 6011
,( 4, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(24,24),(14,17)), 0, 12) -- 6012
,( 4, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(26,26),(16,19)), 0, 12) -- 6013
,( 4, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 6014
,( 4, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 6015
,( 4, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 6016
,( 4, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 6017
,( 4, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 6018
,( 4, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 6019
,( 4, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 6020
,( 4, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 6021
,( 4, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 6022
,( 4, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(22,23),(10,13)), 0, 11) -- 6023
,( 4, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(24,25),(12,15)), 0, 11) -- 6024
,( 4, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(26,27),(14,17)), 0, 11) -- 6025
,( 4, E,0,0,((24,27),(22,22),( 1, 1),(18,19),(22,23),(12,13)), 0, 11) -- 6026
,( 4, E,0,0,((26,29),(24,24),( 3, 3),(20,21),(24,25),(14,15)), 0, 11) -- 6027
,( 4, E,0,0,((28,31),(26,26),( 5, 5),(22,23),(26,27),(16,17)), 0, 11) -- 6028
,( 4, E,0,0,((30,33),(28,28),( 7, 7),(24,25),(28,29),(18,19)), 0, 11) -- 6029
,( 4, E,0,0,((22,25),(18,19),( 0, 1),(18,19),(22,22),(14,17)), 0, 11) -- 6030
,( 4, E,0,0,((24,27),(20,21),( 2, 3),(20,21),(24,24),(16,19)), 0, 11) -- 6031
,( 4, E,0,0,((26,29),(22,23),( 4, 5),(22,23),(26,26),(18,21)), 0, 11) -- 6032
,( 4, E,0,0,((28,31),(24,25),( 6, 7),(24,25),(28,28),(20,23)), 0, 11) -- 6033
,( 4, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(10,13)), 0, 10) -- 6034
,( 4, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(12,15)), 0, 10) -- 6035
,( 4, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(14,17)), 0, 10) -- 6036
,( 4, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(16,19)), 0, 10) -- 6037
,( 4, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(21,21),(10,13)), 0, 10) -- 6038
,( 4, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(23,23),(12,15)), 0, 10) -- 6039
,( 4, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(25,25),(14,17)), 0, 10) -- 6040
,( 4, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(27,27),(16,19)), 0, 10) -- 6041
,( 4, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 6042
,( 4, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 6043
,( 4, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 6044
,( 4, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 6045
,( 4, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 6, 9)), 0, 10) -- 6046
,( 4, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),( 8,11)), 0, 10) -- 6047
,( 4, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(10,13)), 0, 10) -- 6048
,( 4, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(12,15)), 0, 10) -- 6049
,( 4, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(20,20),( 8,11)), 0, 10) -- 6050
,( 4, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(22,22),(10,13)), 0, 10) -- 6051
,( 4, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(24,24),(12,15)), 0, 10) -- 6052
,( 4, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(26,26),(14,17)), 0, 10) -- 6053
,( 4, E,0,0,((22,23),(20,20),( 0, 1),(18,19),(22,23),(14,17)), 0, 10) -- 6054
,( 4, E,0,0,((24,25),(22,22),( 2, 3),(20,21),(24,25),(16,19)), 0, 10) -- 6055
,( 4, E,0,0,((26,27),(24,24),( 4, 5),(22,23),(26,27),(18,21)), 0, 10) -- 6056
,( 4, E,0,0,((28,29),(26,26),( 6, 7),(24,25),(28,29),(20,23)), 0, 10) -- 6057
,( 4, E,0,0,((24,27),(20,21),( 0, 1),(17,17),(16,16),( 4, 7)), 0, 10) -- 6058
,( 4, E,0,0,((26,29),(22,23),( 2, 3),(19,19),(18,18),( 6, 9)), 0, 10) -- 6059
,( 4, E,0,0,((28,31),(24,25),( 4, 5),(21,21),(20,20),( 8,11)), 0, 10) -- 6060
,( 4, E,0,0,((30,33),(26,27),( 6, 7),(23,23),(22,22),(10,13)), 0, 10) -- 6061
,( 4, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(18,19),( 4, 7)), 0, 10) -- 6062
,( 4, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(20,21),( 6, 9)), 0, 10) -- 6063
,( 4, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(22,23),( 8,11)), 0, 10) -- 6064
,( 4, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(24,25),(10,13)), 0, 10) -- 6065
,( 4, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(12,15)), 0, 10) -- 6066
,( 4, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(14,17)), 0, 10) -- 6067
,( 4, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(16,19)), 0, 10) -- 6068
,( 4, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(18,21)), 0, 10) -- 6069
,( 4, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),( 4, 7)), 0, 10) -- 6070
,( 4, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),( 6, 9)), 0, 10) -- 6071
,( 4, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),( 8,11)), 0, 10) -- 6072
,( 4, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(10,13)), 0, 10) -- 6073
,( 4, E,0,0,((24,27),(22,22),( 0, 1),(18,19),(22,23),( 8,11)), 0, 10) -- 6074
,( 4, E,0,0,((26,29),(24,24),( 2, 3),(20,21),(24,25),(10,13)), 0, 10) -- 6075
,( 4, E,0,0,((28,31),(26,26),( 4, 5),(22,23),(26,27),(12,15)), 0, 10) -- 6076
,( 4, E,0,0,((30,33),(28,28),( 6, 7),(24,25),(28,29),(14,17)), 0, 10) -- 6077
,( 4, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(24,24),(16,19)), 0, 10) -- 6078
,( 4, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(26,26),(18,21)), 0, 10) -- 6079
,( 4, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(28,28),(20,23)), 0, 10) -- 6080
,( 4, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(30,30),(22,23)), 0, 10) -- 6081
,( 4, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(99,99),( 8,11)), 0, 10) -- 6082
,( 4, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(99,99),(10,13)), 0, 10) -- 6083
,( 4, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(99,99),(12,15)), 0, 10) -- 6084
,( 4, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(99,99),(14,17)), 0, 10) -- 6085
,( 4, E,0,0,((18,21),(18,19),( 0, 1),(20,20),(24,25),(14,17)), 0,  9) -- 6086
,( 4, E,0,0,((20,23),(20,21),( 2, 3),(22,22),(26,27),(16,19)), 0,  9) -- 6087
,( 4, E,0,0,((22,25),(22,23),( 4, 5),(24,24),(28,29),(18,21)), 0,  9) -- 6088
,( 4, E,0,0,((24,27),(24,25),( 6, 7),(26,26),(30,31),(20,23)), 0,  9) -- 6089
,( 4, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 6090
,( 4, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 6091
,( 4, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 6092
,( 4, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 6093
,( 4, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(22,23),(10,13)), 0,  9) -- 6094
,( 4, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(24,25),(12,15)), 0,  9) -- 6095
,( 4, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(26,27),(14,17)), 0,  9) -- 6096
,( 4, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(28,29),(16,19)), 0,  9) -- 6097
,( 4, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 6098
,( 4, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 6099
,( 4, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 6100
,( 4, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 6101
,( 4, E,0,0,((16,19),(16,17),( 0, 1),(18,19),(24,25),(12,15)), 0,  9) -- 6102
,( 4, E,0,0,((18,21),(18,19),( 2, 3),(20,21),(26,27),(14,17)), 0,  9) -- 6103
,( 4, E,0,0,((20,23),(20,21),( 4, 5),(22,23),(28,29),(16,19)), 0,  9) -- 6104
,( 4, E,0,0,((22,25),(22,23),( 6, 7),(24,25),(30,31),(18,21)), 0,  9) -- 6105
,( 4, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(24,25),(14,17)), 0,  9) -- 6106
,( 4, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(26,27),(16,19)), 0,  9) -- 6107
,( 4, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(28,29),(18,21)), 0,  9) -- 6108
,( 4, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(30,31),(20,23)), 0,  9) -- 6109
,( 4, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),( 6, 9)), 0,  9) -- 6110
,( 4, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),( 8,11)), 0,  9) -- 6111
,( 4, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(10,13)), 0,  9) -- 6112
,( 4, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(12,15)), 0,  9) -- 6113
,( 4, E,0,0,((20,23),(18,19),( 0, 0),(18,18),(20,21),( 6, 9)), 0,  9) -- 6114
,( 4, E,0,0,((22,25),(20,21),( 2, 2),(20,20),(22,23),( 8,11)), 0,  9) -- 6115
,( 4, E,0,0,((24,27),(22,23),( 4, 4),(22,22),(24,25),(10,13)), 0,  9) -- 6116
,( 4, E,0,0,((26,29),(24,25),( 6, 6),(24,24),(26,27),(12,15)), 0,  9) -- 6117
,( 4, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(22,23),(12,15)), 0,  9) -- 6118
,( 4, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(24,25),(14,17)), 0,  9) -- 6119
,( 4, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(26,27),(16,19)), 0,  9) -- 6120
,( 4, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(28,29),(18,21)), 0,  9) -- 6121
,( 4, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 6122
,( 4, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 6123
,( 4, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 6124
,( 4, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 6125
,( 4, E,0,0,((20,23),(20,20),( 1, 1),(20,21),(24,25),(14,17)), 0,  9) -- 6126
,( 4, E,0,0,((22,25),(22,22),( 3, 3),(22,23),(26,27),(16,19)), 0,  9) -- 6127
,( 4, E,0,0,((24,27),(24,24),( 5, 5),(24,25),(28,29),(18,21)), 0,  9) -- 6128
,( 4, E,0,0,((26,29),(26,26),( 7, 7),(26,27),(30,31),(20,23)), 0,  9) -- 6129
,( 4, E,0,0,((20,23),(18,19),( 0, 1),(20,21),(24,25),(10,13)), 0,  9) -- 6130
,( 4, E,0,0,((22,25),(20,21),( 2, 3),(22,23),(26,27),(12,15)), 0,  9) -- 6131
,( 4, E,0,0,((24,27),(22,23),( 4, 5),(24,25),(28,29),(14,17)), 0,  9) -- 6132
,( 4, E,0,0,((26,29),(24,25),( 6, 7),(26,27),(30,31),(16,19)), 0,  9) -- 6133
,( 4, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(20,21),(10,13)), 0,  9) -- 6134
,( 4, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(22,23),(12,15)), 0,  9) -- 6135
,( 4, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(24,25),(14,17)), 0,  9) -- 6136
,( 4, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(26,27),(16,19)), 0,  9) -- 6137
,( 4, E,0,0,((20,23),(18,19),( 0, 0),(17,17),(20,21),(13,13)), 0,  9) -- 6138
,( 4, E,0,0,((22,25),(20,21),( 2, 2),(19,19),(22,23),(15,15)), 0,  9) -- 6139
,( 4, E,0,0,((24,27),(22,23),( 4, 4),(21,21),(24,25),(17,17)), 0,  9) -- 6140
,( 4, E,0,0,((26,29),(24,25),( 6, 6),(23,23),(26,27),(19,19)), 0,  9) -- 6141
,( 4, E,0,0,((18,21),(18,19),( 1, 1),(20,21),(26,26),(17,17)), 0,  9) -- 6142
,( 4, E,0,0,((20,23),(20,21),( 3, 3),(22,23),(28,28),(19,19)), 0,  9) -- 6143
,( 4, E,0,0,((22,25),(22,23),( 5, 5),(24,25),(30,30),(21,21)), 0,  9) -- 6144
,( 4, E,0,0,((24,27),(24,25),( 7, 7),(26,27),(32,32),(23,23)), 0,  9) -- 6145
,( 4, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(99,99),( 2, 5)), 0,  9) -- 6146
,( 4, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(99,99),( 4, 7)), 0,  9) -- 6147
,( 4, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(99,99),( 6, 9)), 0,  9) -- 6148
,( 4, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(99,99),( 8,11)), 0,  9) -- 6149
,( 4, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(20,23),(99,99)), 0,  8) -- 6150
,( 4, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(22,25),(99,99)), 0,  8) -- 6151
,( 4, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(24,27),(99,99)), 0,  8) -- 6152
,( 4, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(26,29),(99,99)), 0,  8) -- 6153
,( 4, E,0,0,((18,21),(16,19),( 0, 1),(16,19),(16,19),(99,99)), 0,  8) -- 6154
,( 4, E,0,0,((20,23),(18,21),( 2, 3),(18,21),(18,21),(99,99)), 0,  8) -- 6155
,( 4, E,0,0,((22,25),(20,23),( 4, 5),(20,23),(20,23),(99,99)), 0,  8) -- 6156
,( 4, E,0,0,((24,27),(22,25),( 6, 7),(22,25),(22,25),(99,99)), 0,  8) -- 6157
,( 4, E,0,0,((14,17),(14,17),( 0, 1),(18,21),(24,27),(99,99)), 0,  8) -- 6158
,( 4, E,0,0,((16,19),(16,19),( 2, 3),(20,23),(26,29),(99,99)), 0,  8) -- 6159
,( 4, E,0,0,((18,21),(18,21),( 4, 5),(22,25),(28,31),(99,99)), 0,  8) -- 6160
,( 4, E,0,0,((20,23),(20,23),( 6, 7),(24,27),(30,33),(99,99)), 0,  8) -- 6161
,( 4, E,0,0,((18,21),(16,19),( 0, 1),(16,19),(12,15),(99,99)), 0,  7) -- 6162
,( 4, E,0,0,((20,23),(18,21),( 2, 3),(18,21),(14,17),(99,99)), 0,  7) -- 6163
,( 4, E,0,0,((22,25),(20,23),( 4, 5),(20,23),(16,19),(99,99)), 0,  7) -- 6164
,( 4, E,0,0,((24,27),(22,25),( 6, 7),(22,25),(18,21),(99,99)), 0,  7) -- 6165
,( 4, E,0,1,((10,13),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 6166
,( 4, E,0,1,((12,15),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 6167
,( 4, E,0,1,((14,17),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 6168
,( 4, E,0,1,((16,19),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 6169
,( 4, E,0,1,((14,17),(16,19),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 6170
,( 4, E,0,1,((16,19),(18,21),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 6171
,( 4, E,0,1,((18,21),(20,23),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 6172
,( 4, E,0,1,((20,23),(22,25),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 6173
,( 4, E,0,1,((18,21),(20,21),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 6174
,( 4, E,0,1,((20,23),(22,23),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 6175
,( 4, E,0,1,((22,25),(24,25),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 6176
,( 4, E,0,1,((24,27),(26,27),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 6177
,( 4, E,0,1,((20,23),(20,23),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 6178
,( 4, E,0,1,((22,25),(22,25),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 6179
,( 4, E,0,1,((24,27),(24,27),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 6180
,( 4, E,0,1,((26,29),(26,29),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 6181
,( 4, E,0,1,((16,19),(16,19),( 0, 0),(12,15),(99,99),(99,99)), 0,  6) -- 6182
,( 4, E,0,1,((18,21),(18,21),( 2, 2),(14,17),(99,99),(99,99)), 0,  6) -- 6183
,( 4, E,0,1,((20,23),(20,23),( 4, 4),(16,19),(99,99),(99,99)), 0,  6) -- 6184
,( 4, E,0,1,((22,25),(22,25),( 6, 6),(18,21),(99,99),(99,99)), 0,  6) -- 6185
,( 4, E,0,1,(( 8,11),(12,15),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 6186
,( 4, E,0,1,((10,13),(14,17),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 6187
,( 4, E,0,1,((12,15),(16,19),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 6188
,( 4, E,0,1,((14,17),(18,21),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 6189
,( 4, E,0,1,((22,25),(22,25),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 6190
,( 4, E,0,1,((24,27),(24,27),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 6191
,( 4, E,0,1,((26,29),(26,29),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 6192
,( 4, E,0,1,((28,31),(28,31),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 6193
,( 4, E,0,1,((24,27),(22,23),( 0, 1),(17,17),(99,99),(99,99)), 0,  5) -- 6194
,( 4, E,0,1,((26,29),(24,25),( 2, 3),(19,19),(99,99),(99,99)), 0,  5) -- 6195
,( 4, E,0,1,((28,31),(26,27),( 4, 5),(21,21),(99,99),(99,99)), 0,  5) -- 6196
,( 4, E,0,1,((30,33),(28,29),( 6, 7),(23,23),(99,99),(99,99)), 0,  5) -- 6197
,( 5, E,0,0,((33,33),(99,99),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 6198
,( 5, E,0,0,((34,34),(99,99),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 6199
,( 5, E,0,0,((35,35),(99,99),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 6200
,( 5, E,0,0,((36,36),(99,99),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 6201
,( 5, E,0,0,((37,37),(99,99),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 6202
,( 5, E,0,0,((38,38),(99,99),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 6203
,( 5, E,0,0,((39,39),(99,99),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 6204
,( 5, E,0,0,((40,40),(99,99),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 6205
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 6206
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 6207
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 6208
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 6209
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 6210
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 6211
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 6212
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 6213
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 30) -- 6214
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 30) -- 6215
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 30) -- 6216
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(18,18),(19,19),(10,10)), 1, 30) -- 6217
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(19,19),(20,20),(11,11)), 1, 30) -- 6218
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(20,20),(21,21),(12,12)), 1, 30) -- 6219
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(21,21),(22,22),(13,13)), 1, 30) -- 6220
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(22,22),(23,23),(14,14)), 1, 30) -- 6221
,( 5, E,0,0,((33,33),(99,99),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 29) -- 6222
,( 5, E,0,0,((34,34),(99,99),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 29) -- 6223
,( 5, E,0,0,((35,35),(99,99),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 29) -- 6224
,( 5, E,0,0,((36,36),(99,99),( 3, 3),(19,19),(19,19),(10,10)), 1, 29) -- 6225
,( 5, E,0,0,((37,37),(99,99),( 4, 4),(20,20),(20,20),(11,11)), 1, 29) -- 6226
,( 5, E,0,0,((38,38),(99,99),( 5, 5),(21,21),(21,21),(12,12)), 1, 29) -- 6227
,( 5, E,0,0,((39,39),(99,99),( 6, 6),(22,22),(22,22),(13,13)), 1, 29) -- 6228
,( 5, E,0,0,((40,40),(99,99),( 7, 7),(23,23),(23,23),(14,14)), 1, 29) -- 6229
,( 5, E,0,0,((33,33),(99,99),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 29) -- 6230
,( 5, E,0,0,((34,34),(99,99),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 29) -- 6231
,( 5, E,0,0,((35,35),(99,99),( 2, 2),(17,17),(18,18),(10,10)), 1, 29) -- 6232
,( 5, E,0,0,((36,36),(99,99),( 3, 3),(18,18),(19,19),(11,11)), 1, 29) -- 6233
,( 5, E,0,0,((37,37),(99,99),( 4, 4),(19,19),(20,20),(12,12)), 1, 29) -- 6234
,( 5, E,0,0,((38,38),(99,99),( 5, 5),(20,20),(21,21),(13,13)), 1, 29) -- 6235
,( 5, E,0,0,((39,39),(99,99),( 6, 6),(21,21),(22,22),(14,14)), 1, 29) -- 6236
,( 5, E,0,0,((40,40),(99,99),( 7, 7),(22,22),(23,23),(15,15)), 1, 29) -- 6237
,( 5, E,0,0,((33,33),(99,99),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 28) -- 6238
,( 5, E,0,0,((34,34),(99,99),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 28) -- 6239
,( 5, E,0,0,((35,35),(99,99),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 28) -- 6240
,( 5, E,0,0,((36,36),(99,99),( 3, 3),(18,18),(19,19),(10,10)), 1, 28) -- 6241
,( 5, E,0,0,((37,37),(99,99),( 4, 4),(19,19),(20,20),(11,11)), 1, 28) -- 6242
,( 5, E,0,0,((38,38),(99,99),( 5, 5),(20,20),(21,21),(12,12)), 1, 28) -- 6243
,( 5, E,0,0,((39,39),(99,99),( 6, 6),(21,21),(22,22),(13,13)), 1, 28) -- 6244
,( 5, E,0,0,((40,40),(99,99),( 7, 7),(22,22),(23,23),(14,14)), 1, 28) -- 6245
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(16,16),(99,99),( 7, 7)), 1, 23) -- 6246
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(17,17),(99,99),( 8, 8)), 1, 23) -- 6247
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(18,18),(99,99),( 9, 9)), 1, 23) -- 6248
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(19,19),(99,99),(10,10)), 1, 23) -- 6249
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(20,20),(99,99),(11,11)), 1, 23) -- 6250
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(21,21),(99,99),(12,12)), 1, 23) -- 6251
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(22,22),(99,99),(13,13)), 1, 23) -- 6252
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(23,23),(99,99),(14,14)), 1, 23) -- 6253
,( 5, E,0,0,((33,33),(99,99),( 0, 0),(15,15),(99,99),( 6, 6)), 1, 22) -- 6254
,( 5, E,0,0,((34,34),(99,99),( 1, 1),(16,16),(99,99),( 7, 7)), 1, 22) -- 6255
,( 5, E,0,0,((35,35),(99,99),( 2, 2),(17,17),(99,99),( 8, 8)), 1, 22) -- 6256
,( 5, E,0,0,((36,36),(99,99),( 3, 3),(18,18),(99,99),( 9, 9)), 1, 22) -- 6257
,( 5, E,0,0,((37,37),(99,99),( 4, 4),(19,19),(99,99),(10,10)), 1, 22) -- 6258
,( 5, E,0,0,((38,38),(99,99),( 5, 5),(20,20),(99,99),(11,11)), 1, 22) -- 6259
,( 5, E,0,0,((39,39),(99,99),( 6, 6),(21,21),(99,99),(12,12)), 1, 22) -- 6260
,( 5, E,0,0,((40,40),(99,99),( 7, 7),(22,22),(99,99),(13,13)), 1, 22) -- 6261
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(16,16),(99,99),( 8, 8)), 1, 21) -- 6262
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(17,17),(99,99),( 9, 9)), 1, 21) -- 6263
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(18,18),(99,99),(10,10)), 1, 21) -- 6264
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(19,19),(99,99),(11,11)), 1, 21) -- 6265
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(20,20),(99,99),(12,12)), 1, 21) -- 6266
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(21,21),(99,99),(13,13)), 1, 21) -- 6267
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(22,22),(99,99),(14,14)), 1, 21) -- 6268
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(23,23),(99,99),(15,15)), 1, 21) -- 6269
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(15,15),(99,99),( 7, 7)), 1, 20) -- 6270
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(16,16),(99,99),( 8, 8)), 1, 20) -- 6271
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(17,17),(99,99),( 9, 9)), 1, 20) -- 6272
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(18,18),(99,99),(10,10)), 1, 20) -- 6273
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(19,19),(99,99),(11,11)), 1, 20) -- 6274
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(20,20),(99,99),(12,12)), 1, 20) -- 6275
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(21,21),(99,99),(13,13)), 1, 20) -- 6276
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(22,22),(99,99),(14,14)), 1, 20) -- 6277
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(15,15),(99,99),( 6, 6)), 1, 19) -- 6278
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(16,16),(99,99),( 7, 7)), 1, 19) -- 6279
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(17,17),(99,99),( 8, 8)), 1, 19) -- 6280
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(18,18),(99,99),( 9, 9)), 1, 19) -- 6281
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(19,19),(99,99),(10,10)), 1, 19) -- 6282
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(20,20),(99,99),(11,11)), 1, 19) -- 6283
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(21,21),(99,99),(12,12)), 1, 19) -- 6284
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(22,22),(99,99),(13,13)), 1, 19) -- 6285
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(15,15),(99,99),( 8, 8)), 1, 18) -- 6286
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(16,16),(99,99),( 9, 9)), 1, 18) -- 6287
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(17,17),(99,99),(10,10)), 1, 18) -- 6288
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(18,18),(99,99),(11,11)), 1, 18) -- 6289
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(19,19),(99,99),(12,12)), 1, 18) -- 6290
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(20,20),(99,99),(13,13)), 1, 18) -- 6291
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(21,21),(99,99),(14,14)), 1, 18) -- 6292
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(22,22),(99,99),(15,15)), 1, 18) -- 6293
,( 5, E,0,0,((35,35),(99,99),( 0, 0),(15,15),(99,99),( 6, 6)), 1, 18) -- 6294
,( 5, E,0,0,((36,36),(99,99),( 1, 1),(16,16),(99,99),( 7, 7)), 1, 18) -- 6295
,( 5, E,0,0,((37,37),(99,99),( 2, 2),(17,17),(99,99),( 8, 8)), 1, 18) -- 6296
,( 5, E,0,0,((38,38),(99,99),( 3, 3),(18,18),(99,99),( 9, 9)), 1, 18) -- 6297
,( 5, E,0,0,((39,39),(99,99),( 4, 4),(19,19),(99,99),(10,10)), 1, 18) -- 6298
,( 5, E,0,0,((40,40),(99,99),( 5, 5),(20,20),(99,99),(11,11)), 1, 18) -- 6299
,( 5, E,0,0,((41,41),(99,99),( 6, 6),(21,21),(99,99),(12,12)), 1, 18) -- 6300
,( 5, E,0,0,((42,42),(99,99),( 7, 7),(22,22),(99,99),(13,13)), 1, 18) -- 6301
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(15,15),(99,99),( 5, 5)), 1, 18) -- 6302
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(16,16),(99,99),( 6, 6)), 1, 18) -- 6303
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(17,17),(99,99),( 7, 7)), 1, 18) -- 6304
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(18,18),(99,99),( 8, 8)), 1, 18) -- 6305
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(19,19),(99,99),( 9, 9)), 1, 18) -- 6306
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(20,20),(99,99),(10,10)), 1, 18) -- 6307
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(21,21),(99,99),(11,11)), 1, 18) -- 6308
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(22,22),(99,99),(12,12)), 1, 18) -- 6309
,( 5, E,0,0,((35,35),(99,99),( 0, 0),(15,15),(99,99),( 7, 7)), 1, 17) -- 6310
,( 5, E,0,0,((36,36),(99,99),( 1, 1),(16,16),(99,99),( 8, 8)), 1, 17) -- 6311
,( 5, E,0,0,((37,37),(99,99),( 2, 2),(17,17),(99,99),( 9, 9)), 1, 17) -- 6312
,( 5, E,0,0,((38,38),(99,99),( 3, 3),(18,18),(99,99),(10,10)), 1, 17) -- 6313
,( 5, E,0,0,((39,39),(99,99),( 4, 4),(19,19),(99,99),(11,11)), 1, 17) -- 6314
,( 5, E,0,0,((40,40),(99,99),( 5, 5),(20,20),(99,99),(12,12)), 1, 17) -- 6315
,( 5, E,0,0,((41,41),(99,99),( 6, 6),(21,21),(99,99),(13,13)), 1, 17) -- 6316
,( 5, E,0,0,((42,42),(99,99),( 7, 7),(22,22),(99,99),(14,14)), 1, 17) -- 6317
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(14,14),(99,99),( 5, 5)), 1, 17) -- 6318
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(15,15),(99,99),( 6, 6)), 1, 17) -- 6319
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(16,16),(99,99),( 7, 7)), 1, 17) -- 6320
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(17,17),(99,99),( 8, 8)), 1, 17) -- 6321
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(18,18),(99,99),( 9, 9)), 1, 17) -- 6322
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(19,19),(99,99),(10,10)), 1, 17) -- 6323
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(20,20),(99,99),(11,11)), 1, 17) -- 6324
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(21,21),(99,99),(12,12)), 1, 17) -- 6325
,( 5, E,0,0,((34,34),(99,99),( 0, 0),(14,14),(99,99),( 6, 6)), 1, 16) -- 6326
,( 5, E,0,0,((35,35),(99,99),( 1, 1),(15,15),(99,99),( 7, 7)), 1, 16) -- 6327
,( 5, E,0,0,((36,36),(99,99),( 2, 2),(16,16),(99,99),( 8, 8)), 1, 16) -- 6328
,( 5, E,0,0,((37,37),(99,99),( 3, 3),(17,17),(99,99),( 9, 9)), 1, 16) -- 6329
,( 5, E,0,0,((38,38),(99,99),( 4, 4),(18,18),(99,99),(10,10)), 1, 16) -- 6330
,( 5, E,0,0,((39,39),(99,99),( 5, 5),(19,19),(99,99),(11,11)), 1, 16) -- 6331
,( 5, E,0,0,((40,40),(99,99),( 6, 6),(20,20),(99,99),(12,12)), 1, 16) -- 6332
,( 5, E,0,0,((41,41),(99,99),( 7, 7),(21,21),(99,99),(13,13)), 1, 16) -- 6333
,( 5, E,0,0,((35,35),(99,99),( 0, 0),(15,15),(99,99),( 5, 5)), 1, 16) -- 6334
,( 5, E,0,0,((36,36),(99,99),( 1, 1),(16,16),(99,99),( 6, 6)), 1, 16) -- 6335
,( 5, E,0,0,((37,37),(99,99),( 2, 2),(17,17),(99,99),( 7, 7)), 1, 16) -- 6336
,( 5, E,0,0,((38,38),(99,99),( 3, 3),(18,18),(99,99),( 8, 8)), 1, 16) -- 6337
,( 5, E,0,0,((39,39),(99,99),( 4, 4),(19,19),(99,99),( 9, 9)), 1, 16) -- 6338
,( 5, E,0,0,((40,40),(99,99),( 5, 5),(20,20),(99,99),(10,10)), 1, 16) -- 6339
,( 5, E,0,0,((41,41),(99,99),( 6, 6),(21,21),(99,99),(11,11)), 1, 16) -- 6340
,( 5, E,0,0,((42,42),(99,99),( 7, 7),(22,22),(99,99),(12,12)), 1, 16) -- 6341
,( 5, E,0,0,((35,35),(99,99),( 0, 0),(14,14),(99,99),( 6, 6)), 1, 15) -- 6342
,( 5, E,0,0,((36,36),(99,99),( 1, 1),(15,15),(99,99),( 7, 7)), 1, 15) -- 6343
,( 5, E,0,0,((37,37),(99,99),( 2, 2),(16,16),(99,99),( 8, 8)), 1, 15) -- 6344
,( 5, E,0,0,((38,38),(99,99),( 3, 3),(17,17),(99,99),( 9, 9)), 1, 15) -- 6345
,( 5, E,0,0,((39,39),(99,99),( 4, 4),(18,18),(99,99),(10,10)), 1, 15) -- 6346
,( 5, E,0,0,((40,40),(99,99),( 5, 5),(19,19),(99,99),(11,11)), 1, 15) -- 6347
,( 5, E,0,0,((41,41),(99,99),( 6, 6),(20,20),(99,99),(12,12)), 1, 15) -- 6348
,( 5, E,0,0,((42,42),(99,99),( 7, 7),(21,21),(99,99),(13,13)), 1, 15) -- 6349
,( 5, E,0,0,((35,35),(99,99),( 0, 0),(14,14),(99,99),( 5, 5)), 1, 15) -- 6350
,( 5, E,0,0,((36,36),(99,99),( 1, 1),(15,15),(99,99),( 6, 6)), 1, 15) -- 6351
,( 5, E,0,0,((37,37),(99,99),( 2, 2),(16,16),(99,99),( 7, 7)), 1, 15) -- 6352
,( 5, E,0,0,((38,38),(99,99),( 3, 3),(17,17),(99,99),( 8, 8)), 1, 15) -- 6353
,( 5, E,0,0,((39,39),(99,99),( 4, 4),(18,18),(99,99),( 9, 9)), 1, 15) -- 6354
,( 5, E,0,0,((40,40),(99,99),( 5, 5),(19,19),(99,99),(10,10)), 1, 15) -- 6355
,( 5, E,0,0,((41,41),(99,99),( 6, 6),(20,20),(99,99),(11,11)), 1, 15) -- 6356
,( 5, E,0,0,((42,42),(99,99),( 7, 7),(21,21),(99,99),(12,12)), 1, 15) -- 6357
,( 5, E,0,0,((34,37),(99,99),( 0, 1),(14,15),(14,14),( 4, 7)), 1, 14) -- 6358
,( 5, E,0,0,((36,39),(99,99),( 2, 3),(16,17),(16,16),( 6, 9)), 1, 14) -- 6359
,( 5, E,0,0,((38,41),(99,99),( 4, 5),(18,19),(18,18),( 8,11)), 1, 14) -- 6360
,( 5, E,0,0,((40,43),(99,99),( 6, 7),(20,21),(20,20),(10,13)), 1, 14) -- 6361
,( 5, E,0,0,((38,38),(99,99),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 6362
,( 5, E,0,0,((40,40),(99,99),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 6363
,( 5, E,0,0,((42,42),(99,99),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 6364
,( 5, E,0,0,((44,44),(99,99),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 6365
,( 5, E,0,0,((36,39),(99,99),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 6366
,( 5, E,0,0,((38,41),(99,99),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 6367
,( 5, E,0,0,((40,43),(99,99),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 6368
,( 5, E,0,0,((42,45),(99,99),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 6369
,( 5, E,0,0,((36,39),(99,99),( 1, 1),(15,15),(14,14),( 6, 9)), 1, 14) -- 6370
,( 5, E,0,0,((38,41),(99,99),( 3, 3),(17,17),(16,16),( 8,11)), 1, 14) -- 6371
,( 5, E,0,0,((40,43),(99,99),( 5, 5),(19,19),(18,18),(10,13)), 1, 14) -- 6372
,( 5, E,0,0,((42,45),(99,99),( 7, 7),(21,21),(20,20),(12,15)), 1, 14) -- 6373
,( 5, E,0,0,((38,41),(99,99),( 0, 1),(15,15),(14,15),( 4, 7)), 1, 13) -- 6374
,( 5, E,0,0,((40,43),(99,99),( 2, 3),(17,17),(16,17),( 6, 9)), 1, 13) -- 6375
,( 5, E,0,0,((42,45),(99,99),( 4, 5),(19,19),(18,19),( 8,11)), 1, 13) -- 6376
,( 5, E,0,0,((44,47),(99,99),( 6, 7),(21,21),(20,21),(10,13)), 1, 13) -- 6377
,( 5, E,0,0,((39,39),(99,99),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 13) -- 6378
,( 5, E,0,0,((41,41),(99,99),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 13) -- 6379
,( 5, E,0,0,((43,43),(99,99),( 5, 5),(20,20),(18,19),( 8,11)), 1, 13) -- 6380
,( 5, E,0,0,((45,45),(99,99),( 7, 7),(22,22),(20,21),(10,13)), 1, 13) -- 6381
,( 5, E,0,0,((38,41),(99,99),( 0, 1),(14,15),(12,13),( 4, 7)), 1, 12) -- 6382
,( 5, E,0,0,((40,43),(99,99),( 2, 3),(16,17),(14,15),( 6, 9)), 1, 12) -- 6383
,( 5, E,0,0,((42,45),(99,99),( 4, 5),(18,19),(16,17),( 8,11)), 1, 12) -- 6384
,( 5, E,0,0,((44,47),(99,99),( 6, 7),(20,21),(18,19),(10,13)), 1, 12) -- 6385
,( 5, E,0,0,((40,41),(99,99),( 0, 1),(14,15),(12,13),( 0, 3)), 1, 12) -- 6386
,( 5, E,0,0,((42,43),(99,99),( 2, 3),(16,17),(14,15),( 2, 5)), 1, 12) -- 6387
,( 5, E,0,0,((44,45),(99,99),( 4, 5),(18,19),(16,17),( 4, 7)), 1, 12) -- 6388
,( 5, E,0,0,((46,47),(99,99),( 6, 7),(20,21),(18,19),( 6, 9)), 1, 12) -- 6389
,( 5, E,0,0,((38,41),(99,99),( 0, 0),(13,13),(12,12),( 0, 3)), 1, 12) -- 6390
,( 5, E,0,0,((40,43),(99,99),( 2, 2),(15,15),(14,14),( 2, 5)), 1, 12) -- 6391
,( 5, E,0,0,((42,45),(99,99),( 4, 4),(17,17),(16,16),( 4, 7)), 1, 12) -- 6392
,( 5, E,0,0,((44,47),(99,99),( 6, 6),(19,19),(18,18),( 6, 9)), 1, 12) -- 6393
,( 5, E,0,0,((38,41),(99,99),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 12) -- 6394
,( 5, E,0,0,((40,43),(99,99),( 2, 3),(16,17),(16,17),( 8,11)), 1, 12) -- 6395
,( 5, E,0,0,((42,45),(99,99),( 4, 5),(18,19),(18,19),(10,13)), 1, 12) -- 6396
,( 5, E,0,0,((44,47),(99,99),( 6, 7),(20,21),(20,21),(12,15)), 1, 12) -- 6397
,( 5, E,0,0,((38,41),(99,99),( 0, 0),(13,13),(12,12),( 4, 7)), 1, 11) -- 6398
,( 5, E,0,0,((40,43),(99,99),( 2, 2),(15,15),(14,14),( 6, 9)), 1, 11) -- 6399
,( 5, E,0,0,((42,45),(99,99),( 4, 4),(17,17),(16,16),( 8,11)), 1, 11) -- 6400
,( 5, E,0,0,((44,47),(99,99),( 6, 6),(19,19),(18,18),(10,13)), 1, 11) -- 6401
,( 5, E,0,0,((42,43),(99,99),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 6402
,( 5, E,0,0,((44,45),(99,99),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 6403
,( 5, E,0,0,((46,47),(99,99),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 6404
,( 5, E,0,0,((48,49),(99,99),( 6, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 6405
,( 5, E,0,0,((38,41),(99,99),( 0, 1),(14,15),(14,15),(10,13)), 1, 11) -- 6406
,( 5, E,0,0,((40,43),(99,99),( 2, 3),(16,17),(16,17),(12,15)), 1, 11) -- 6407
,( 5, E,0,0,((42,45),(99,99),( 4, 5),(18,19),(18,19),(14,17)), 1, 11) -- 6408
,( 5, E,0,0,((44,47),(99,99),( 6, 7),(20,21),(20,21),(16,19)), 1, 11) -- 6409
,( 5, E,0,0,((38,41),(99,99),( 0, 1),(14,14),(13,13),( 8,11)), 1, 11) -- 6410
,( 5, E,0,0,((40,43),(99,99),( 2, 3),(16,16),(15,15),(10,13)), 1, 11) -- 6411
,( 5, E,0,0,((42,45),(99,99),( 4, 5),(18,18),(17,17),(12,15)), 1, 11) -- 6412
,( 5, E,0,0,((44,47),(99,99),( 6, 7),(20,20),(19,19),(14,17)), 1, 11) -- 6413
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 6414
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 6415
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,19),(16,17),(10,13)), 1, 10) -- 6416
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,21),(18,19),(12,15)), 1, 10) -- 6417
,( 5, E,0,0,((40,43),(99,99),( 0, 1),(12,13),(11,11),( 4, 7)), 1, 10) -- 6418
,( 5, E,0,0,((42,45),(99,99),( 2, 3),(14,15),(13,13),( 6, 9)), 1, 10) -- 6419
,( 5, E,0,0,((44,47),(99,99),( 4, 5),(16,17),(15,15),( 8,11)), 1, 10) -- 6420
,( 5, E,0,0,((46,49),(99,99),( 6, 7),(18,19),(17,17),(10,13)), 1, 10) -- 6421
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,15),(13,13),(10,13)), 1, 10) -- 6422
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,17),(15,15),(12,15)), 1, 10) -- 6423
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,19),(17,17),(14,17)), 1, 10) -- 6424
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,21),(19,19),(16,19)), 1, 10) -- 6425
,( 5, E,0,0,((40,43),(99,99),( 0, 1),(12,13),(12,13),( 8,11)), 1, 10) -- 6426
,( 5, E,0,0,((42,45),(99,99),( 2, 3),(14,15),(14,15),(10,13)), 1, 10) -- 6427
,( 5, E,0,0,((44,47),(99,99),( 4, 5),(16,17),(16,17),(12,15)), 1, 10) -- 6428
,( 5, E,0,0,((46,49),(99,99),( 6, 7),(18,19),(18,19),(14,17)), 1, 10) -- 6429
,( 5, E,0,0,((40,43),(99,99),( 0, 1),(12,13),(11,11),( 0, 3)), 1, 10) -- 6430
,( 5, E,0,0,((42,45),(99,99),( 2, 3),(14,15),(13,13),( 2, 5)), 1, 10) -- 6431
,( 5, E,0,0,((44,47),(99,99),( 4, 5),(16,17),(15,15),( 4, 7)), 1, 10) -- 6432
,( 5, E,0,0,((46,49),(99,99),( 6, 7),(18,19),(17,17),( 6, 9)), 1, 10) -- 6433
,( 5, E,0,0,((40,43),(99,99),( 0, 1),(14,15),(14,15),(14,17)), 1, 10) -- 6434
,( 5, E,0,0,((42,45),(99,99),( 2, 3),(16,17),(16,17),(16,19)), 1, 10) -- 6435
,( 5, E,0,0,((44,47),(99,99),( 4, 5),(18,19),(18,19),(18,21)), 1, 10) -- 6436
,( 5, E,0,0,((46,49),(99,99),( 6, 7),(20,21),(20,21),(20,23)), 1, 10) -- 6437
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(13,13),(99,99),(12,15)), 1, 10) -- 6438
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(15,15),(99,99),(14,17)), 1, 10) -- 6439
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(17,17),(99,99),(16,19)), 1, 10) -- 6440
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(19,19),(99,99),(18,21)), 1, 10) -- 6441
,( 5, E,0,0,((44,45),(99,99),( 0, 1),(13,13),(99,99),( 6, 9)), 1, 10) -- 6442
,( 5, E,0,0,((46,47),(99,99),( 2, 3),(15,15),(99,99),( 8,11)), 1, 10) -- 6443
,( 5, E,0,0,((48,49),(99,99),( 4, 5),(17,17),(99,99),(10,13)), 1, 10) -- 6444
,( 5, E,0,0,((50,51),(99,99),( 6, 7),(19,19),(99,99),(12,15)), 1, 10) -- 6445
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 6446
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 6447
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 6448
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 6449
,( 5, E,0,0,((44,47),(30,31),( 0, 1),(12,13),(99,99),( 4, 7)), 1,  9) -- 6450
,( 5, E,0,0,((46,49),(32,33),( 2, 3),(14,15),(99,99),( 6, 9)), 1,  9) -- 6451
,( 5, E,0,0,((48,51),(34,35),( 4, 5),(16,17),(99,99),( 8,11)), 1,  9) -- 6452
,( 5, E,0,0,((50,53),(36,37),( 6, 7),(18,19),(99,99),(10,13)), 1,  9) -- 6453
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(12,13),(12,13),(10,13)), 1,  9) -- 6454
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(14,15),(14,15),(12,15)), 1,  9) -- 6455
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(16,17),(16,17),(14,17)), 1,  9) -- 6456
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(18,19),(18,19),(16,19)), 1,  9) -- 6457
,( 5, E,0,0,((40,43),(99,99),( 0, 0),(13,13),(13,13),(14,17)), 1,  9) -- 6458
,( 5, E,0,0,((42,45),(99,99),( 2, 2),(15,15),(15,15),(16,19)), 1,  9) -- 6459
,( 5, E,0,0,((44,47),(99,99),( 4, 4),(17,17),(17,17),(18,21)), 1,  9) -- 6460
,( 5, E,0,0,((46,49),(99,99),( 6, 6),(19,19),(19,19),(20,23)), 1,  9) -- 6461
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,14),(11,11),( 2, 5)), 1,  9) -- 6462
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,16),(13,13),( 4, 7)), 1,  9) -- 6463
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,18),(15,15),( 6, 9)), 1,  9) -- 6464
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,20),(17,17),( 8,11)), 1,  9) -- 6465
,( 5, E,0,0,((40,43),(99,99),( 0, 0),(14,14),(12,13),(10,13)), 1,  9) -- 6466
,( 5, E,0,0,((42,45),(99,99),( 2, 2),(16,16),(14,15),(12,15)), 1,  9) -- 6467
,( 5, E,0,0,((44,47),(99,99),( 4, 4),(18,18),(16,17),(14,17)), 1,  9) -- 6468
,( 5, E,0,0,((46,49),(99,99),( 6, 6),(20,20),(18,19),(16,19)), 1,  9) -- 6469
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 6470
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 6471
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(16,17),(14,15),(10,13)), 1,  9) -- 6472
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(18,19),(16,17),(12,15)), 1,  9) -- 6473
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,14),(14,14),(16,19)), 1,  9) -- 6474
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,16),(16,16),(18,21)), 1,  9) -- 6475
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,18),(18,18),(20,23)), 1,  9) -- 6476
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,20),(20,20),(22,23)), 1,  9) -- 6477
,( 5, E,0,0,((38,41),(99,99),( 0, 0),(13,13),(12,13),(12,15)), 1,  9) -- 6478
,( 5, E,0,0,((40,43),(99,99),( 2, 2),(15,15),(14,15),(14,17)), 1,  9) -- 6479
,( 5, E,0,0,((42,45),(99,99),( 4, 4),(17,17),(16,17),(16,19)), 1,  9) -- 6480
,( 5, E,0,0,((44,47),(99,99),( 6, 6),(19,19),(18,19),(18,21)), 1,  9) -- 6481
,( 5, E,0,0,((44,47),(99,99),( 1, 1),(14,15),(12,13),(12,15)), 1,  9) -- 6482
,( 5, E,0,0,((46,49),(99,99),( 3, 3),(16,17),(14,15),(14,17)), 1,  9) -- 6483
,( 5, E,0,0,((48,51),(99,99),( 5, 5),(18,19),(16,17),(16,19)), 1,  9) -- 6484
,( 5, E,0,0,((50,53),(99,99),( 7, 7),(20,21),(18,19),(18,21)), 1,  9) -- 6485
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(13,13),(12,12),( 6, 9)), 1,  9) -- 6486
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(15,15),(14,14),( 8,11)), 1,  9) -- 6487
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(17,17),(16,16),(10,13)), 1,  9) -- 6488
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(19,19),(18,18),(12,15)), 1,  9) -- 6489
,( 5, E,0,0,((44,47),(99,99),( 0, 0),(12,13),( 9, 9),( 8, 8)), 1,  9) -- 6490
,( 5, E,0,0,((46,49),(99,99),( 2, 2),(14,15),(11,11),(10,10)), 1,  9) -- 6491
,( 5, E,0,0,((48,51),(99,99),( 4, 4),(16,17),(13,13),(12,12)), 1,  9) -- 6492
,( 5, E,0,0,((50,53),(99,99),( 6, 6),(18,19),(15,15),(14,14)), 1,  9) -- 6493
,( 5, E,0,0,((40,43),(99,99),( 0, 1),(14,15),(16,17),(99,99)), 1,  9) -- 6494
,( 5, E,0,0,((42,45),(99,99),( 2, 3),(16,17),(18,19),(99,99)), 1,  9) -- 6495
,( 5, E,0,0,((44,47),(99,99),( 4, 5),(18,19),(20,21),(99,99)), 1,  9) -- 6496
,( 5, E,0,0,((46,49),(99,99),( 6, 7),(20,21),(22,23),(99,99)), 1,  9) -- 6497
,( 5, E,0,0,((40,43),(99,99),( 0, 0),(13,13),(14,15),(99,99)), 1,  9) -- 6498
,( 5, E,0,0,((42,45),(99,99),( 2, 2),(15,15),(16,17),(99,99)), 1,  9) -- 6499
,( 5, E,0,0,((44,47),(99,99),( 4, 4),(17,17),(18,19),(99,99)), 1,  9) -- 6500
,( 5, E,0,0,((46,49),(99,99),( 6, 6),(19,19),(20,21),(99,99)), 1,  9) -- 6501
,( 5, E,0,0,((44,47),(30,31),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 6502
,( 5, E,0,0,((46,49),(32,33),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 6503
,( 5, E,0,0,((48,51),(34,35),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 6504
,( 5, E,0,0,((50,53),(36,37),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 6505
,( 5, E,0,0,((46,49),(30,33),( 0, 1),(10,13),(10,13),(99,99)), 1,  8) -- 6506
,( 5, E,0,0,((48,51),(32,35),( 2, 3),(12,15),(12,15),(99,99)), 1,  8) -- 6507
,( 5, E,0,0,((50,53),(34,37),( 4, 5),(14,17),(14,17),(99,99)), 1,  8) -- 6508
,( 5, E,0,0,((52,55),(36,39),( 6, 7),(16,19),(16,19),(99,99)), 1,  8) -- 6509
,( 5, E,0,0,((48,51),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 6510
,( 5, E,0,0,((50,53),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 6511
,( 5, E,0,0,((52,55),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 6512
,( 5, E,0,0,((54,57),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 6513
,( 5, E,0,0,((42,45),(99,99),( 0, 1),(14,17),(16,19),(99,99)), 1,  8) -- 6514
,( 5, E,0,0,((44,47),(99,99),( 2, 3),(16,19),(18,21),(99,99)), 1,  8) -- 6515
,( 5, E,0,0,((46,49),(99,99),( 4, 5),(18,21),(20,23),(99,99)), 1,  8) -- 6516
,( 5, E,0,0,((48,51),(99,99),( 6, 7),(20,23),(22,25),(99,99)), 1,  8) -- 6517
,( 5, E,0,0,((44,47),(99,99),( 0, 1),(12,15),(18,21),(99,99)), 1,  8) -- 6518
,( 5, E,0,0,((46,49),(99,99),( 2, 3),(14,17),(20,23),(99,99)), 1,  8) -- 6519
,( 5, E,0,0,((48,51),(99,99),( 4, 5),(16,19),(22,25),(99,99)), 1,  8) -- 6520
,( 5, E,0,0,((50,53),(99,99),( 6, 7),(18,21),(24,27),(99,99)), 1,  8) -- 6521
,( 5, E,0,1,((50,53),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 6522
,( 5, E,0,1,((52,55),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 6523
,( 5, E,0,1,((54,57),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 6524
,( 5, E,0,1,((56,59),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 6525
,( 5, E,0,1,((50,53),(32,35),( 0, 1),( 8,11),(99,99),(99,99)), 1,  7) -- 6526
,( 5, E,0,1,((52,55),(34,37),( 2, 3),(10,13),(99,99),(99,99)), 1,  7) -- 6527
,( 5, E,0,1,((54,57),(36,39),( 4, 5),(12,15),(99,99),(99,99)), 1,  7) -- 6528
,( 5, E,0,1,((56,59),(38,41),( 6, 7),(14,17),(99,99),(99,99)), 1,  7) -- 6529
,( 5, E,0,1,((46,49),(99,99),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 6530
,( 5, E,0,1,((48,51),(99,99),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 6531
,( 5, E,0,1,((50,53),(99,99),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 6532
,( 5, E,0,1,((52,55),(99,99),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 6533
,( 5, E,0,1,((42,45),(99,99),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 6534
,( 5, E,0,1,((44,47),(99,99),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 6535
,( 5, E,0,1,((46,49),(99,99),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 6536
,( 5, E,0,1,((48,51),(99,99),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 6537
,( 5, E,0,1,((46,49),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 1,  7) -- 6538
,( 5, E,0,1,((48,51),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 1,  7) -- 6539
,( 5, E,0,1,((50,53),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 1,  7) -- 6540
,( 5, E,0,1,((52,55),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 1,  7) -- 6541
,( 5, E,0,1,((42,45),(99,99),( 0, 1),(16,17),(99,99),(99,99)), 1,  7) -- 6542
,( 5, E,0,1,((44,47),(99,99),( 2, 3),(18,19),(99,99),(99,99)), 1,  7) -- 6543
,( 5, E,0,1,((46,49),(99,99),( 4, 5),(20,21),(99,99),(99,99)), 1,  7) -- 6544
,( 5, E,0,1,((48,51),(99,99),( 6, 7),(22,23),(99,99),(99,99)), 1,  7) -- 6545
,( 5, E,0,1,((54,57),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  6) -- 6546
,( 5, E,0,1,((56,59),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  6) -- 6547
,( 5, E,0,1,((58,61),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  6) -- 6548
,( 5, E,0,1,((60,63),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  6) -- 6549
,( 5, E,0,1,((50,53),(30,33),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 6550
,( 5, E,0,1,((52,55),(32,35),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 6551
,( 5, E,0,1,((54,57),(34,37),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 6552
,( 5, E,0,1,((56,59),(36,39),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 6553
,( 5, E,0,1,((42,45),(99,99),( 0, 1),(18,21),(99,99),(99,99)), 1,  6) -- 6554
,( 5, E,0,1,((44,47),(99,99),( 2, 3),(20,23),(99,99),(99,99)), 1,  6) -- 6555
,( 5, E,0,1,((46,49),(99,99),( 4, 5),(22,25),(99,99),(99,99)), 1,  6) -- 6556
,( 5, E,0,1,((48,51),(99,99),( 6, 7),(24,27),(99,99),(99,99)), 1,  6) -- 6557
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 6558
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 6559
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 6560
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 6561
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 6562
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 6563
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 6564
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 6565
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 6566
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 6567
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 6568
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 6569
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 6570
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 6571
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 6572
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 6573
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 6574
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 6575
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 6576
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 6577
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 6578
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 6579
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 6580
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 6581
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 30) -- 6582
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 30) -- 6583
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(18,18),(19,19),(10,10)), 0, 30) -- 6584
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(19,19),(20,20),(11,11)), 0, 30) -- 6585
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(20,20),(21,21),(12,12)), 0, 30) -- 6586
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(21,21),(22,22),(13,13)), 0, 30) -- 6587
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(22,22),(23,23),(14,14)), 0, 30) -- 6588
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(23,23),(24,24),(15,15)), 0, 30) -- 6589
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 30) -- 6590
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(17,17),(17,17),(10,10)), 0, 30) -- 6591
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(18,18),(18,18),(11,11)), 0, 30) -- 6592
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(19,19),(19,19),(12,12)), 0, 30) -- 6593
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(20,20),(20,20),(13,13)), 0, 30) -- 6594
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(21,21),(21,21),(14,14)), 0, 30) -- 6595
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(22,22),(22,22),(15,15)), 0, 30) -- 6596
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(23,23),(23,23),(16,16)), 0, 30) -- 6597
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 29) -- 6598
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 29) -- 6599
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(17,17),(18,18),(10,10)), 0, 29) -- 6600
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(18,18),(19,19),(11,11)), 0, 29) -- 6601
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(19,19),(20,20),(12,12)), 0, 29) -- 6602
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(20,20),(21,21),(13,13)), 0, 29) -- 6603
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(21,21),(22,22),(14,14)), 0, 29) -- 6604
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(22,22),(23,23),(15,15)), 0, 29) -- 6605
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 25) -- 6606
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(17,17),(18,18),(10,10)), 0, 25) -- 6607
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(18,18),(19,19),(11,11)), 0, 25) -- 6608
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(19,19),(20,20),(12,12)), 0, 25) -- 6609
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(20,20),(21,21),(13,13)), 0, 25) -- 6610
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(21,21),(22,22),(14,14)), 0, 25) -- 6611
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(22,22),(23,23),(15,15)), 0, 25) -- 6612
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(23,23),(24,24),(16,16)), 0, 25) -- 6613
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 25) -- 6614
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(16,16),(17,17),(10,10)), 0, 25) -- 6615
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(17,17),(18,18),(11,11)), 0, 25) -- 6616
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(18,18),(19,19),(12,12)), 0, 25) -- 6617
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(19,19),(20,20),(13,13)), 0, 25) -- 6618
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(20,20),(21,21),(14,14)), 0, 25) -- 6619
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(21,21),(22,22),(15,15)), 0, 25) -- 6620
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(22,22),(23,23),(16,16)), 0, 25) -- 6621
,( 5, E,0,0,((32,32),(99,99),( 0, 0),(16,16),(17,17),(10,10)), 0, 24) -- 6622
,( 5, E,0,0,((33,33),(99,99),( 1, 1),(17,17),(18,18),(11,11)), 0, 24) -- 6623
,( 5, E,0,0,((34,34),(99,99),( 2, 2),(18,18),(19,19),(12,12)), 0, 24) -- 6624
,( 5, E,0,0,((35,35),(99,99),( 3, 3),(19,19),(20,20),(13,13)), 0, 24) -- 6625
,( 5, E,0,0,((36,36),(99,99),( 4, 4),(20,20),(21,21),(14,14)), 0, 24) -- 6626
,( 5, E,0,0,((37,37),(99,99),( 5, 5),(21,21),(22,22),(15,15)), 0, 24) -- 6627
,( 5, E,0,0,((38,38),(99,99),( 6, 6),(22,22),(23,23),(16,16)), 0, 24) -- 6628
,( 5, E,0,0,((39,39),(99,99),( 7, 7),(23,23),(24,24),(17,17)), 0, 24) -- 6629
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 23) -- 6630
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 23) -- 6631
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(18,18),(19,19),(10,10)), 0, 23) -- 6632
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(19,19),(20,20),(11,11)), 0, 23) -- 6633
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(20,20),(21,21),(12,12)), 0, 23) -- 6634
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(21,21),(22,22),(13,13)), 0, 23) -- 6635
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(22,22),(23,23),(14,14)), 0, 23) -- 6636
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(23,23),(24,24),(15,15)), 0, 23) -- 6637
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(16,16),(17,17),(10,10)), 0, 22) -- 6638
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(17,17),(18,18),(11,11)), 0, 22) -- 6639
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(18,18),(19,19),(12,12)), 0, 22) -- 6640
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(19,19),(20,20),(13,13)), 0, 22) -- 6641
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(20,20),(21,21),(14,14)), 0, 22) -- 6642
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(21,21),(22,22),(15,15)), 0, 22) -- 6643
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(22,22),(23,23),(16,16)), 0, 22) -- 6644
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(23,23),(24,24),(17,17)), 0, 22) -- 6645
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 6646
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 6647
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 6648
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 6649
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 6650
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 6651
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 6652
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 6653
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 20) -- 6654
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(17,17),(18,18),(10,10)), 0, 20) -- 6655
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(18,18),(19,19),(11,11)), 0, 20) -- 6656
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(19,19),(20,20),(12,12)), 0, 20) -- 6657
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(20,20),(21,21),(13,13)), 0, 20) -- 6658
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(21,21),(22,22),(14,14)), 0, 20) -- 6659
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(22,22),(23,23),(15,15)), 0, 20) -- 6660
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(23,23),(24,24),(16,16)), 0, 20) -- 6661
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 6662
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 6663
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 6664
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 6665
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 6666
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 6667
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 6668
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 6669
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 6670
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 6671
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 6672
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 6673
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 6674
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 6675
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 6676
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 6677
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(17,17),(18,18),(11,11)), 0, 19) -- 6678
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(18,18),(19,19),(12,12)), 0, 19) -- 6679
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(19,19),(20,20),(13,13)), 0, 19) -- 6680
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(20,20),(21,21),(14,14)), 0, 19) -- 6681
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(21,21),(22,22),(15,15)), 0, 19) -- 6682
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(22,22),(23,23),(16,16)), 0, 19) -- 6683
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(23,23),(24,24),(17,17)), 0, 19) -- 6684
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(24,24),(25,25),(18,18)), 0, 19) -- 6685
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 6686
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 6687
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 6688
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 6689
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 6690
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 6691
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 6692
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 6693
,( 5, E,0,0,((31,31),(99,99),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 18) -- 6694
,( 5, E,0,0,((32,32),(99,99),( 1, 1),(17,17),(19,19),(10,10)), 0, 18) -- 6695
,( 5, E,0,0,((33,33),(99,99),( 2, 2),(18,18),(20,20),(11,11)), 0, 18) -- 6696
,( 5, E,0,0,((34,34),(99,99),( 3, 3),(19,19),(21,21),(12,12)), 0, 18) -- 6697
,( 5, E,0,0,((35,35),(99,99),( 4, 4),(20,20),(22,22),(13,13)), 0, 18) -- 6698
,( 5, E,0,0,((36,36),(99,99),( 5, 5),(21,21),(23,23),(14,14)), 0, 18) -- 6699
,( 5, E,0,0,((37,37),(99,99),( 6, 6),(22,22),(24,24),(15,15)), 0, 18) -- 6700
,( 5, E,0,0,((38,38),(99,99),( 7, 7),(23,23),(25,25),(16,16)), 0, 18) -- 6701
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(16,16),(18,18),(11,11)), 0, 18) -- 6702
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(17,17),(19,19),(12,12)), 0, 18) -- 6703
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(18,18),(20,20),(13,13)), 0, 18) -- 6704
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(19,19),(21,21),(14,14)), 0, 18) -- 6705
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(20,20),(22,22),(15,15)), 0, 18) -- 6706
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(21,21),(23,23),(16,16)), 0, 18) -- 6707
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(22,22),(24,24),(17,17)), 0, 18) -- 6708
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(23,23),(25,25),(18,18)), 0, 18) -- 6709
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 6710
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 6711
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 6712
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 6713
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 6714
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 6715
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 6716
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 6717
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 6718
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 6719
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 6720
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 6721
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 6722
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 6723
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 6724
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 6725
,( 5, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 6726
,( 5, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 6727
,( 5, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 6728
,( 5, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 6729
,( 5, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 6730
,( 5, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 6731
,( 5, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 6732
,( 5, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 6733
,( 5, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 6734
,( 5, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 6735
,( 5, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 6736
,( 5, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 6737
,( 5, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 6738
,( 5, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 6739
,( 5, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 6740
,( 5, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 6741
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(19,19),(11,11)), 0, 16) -- 6742
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(20,20),(12,12)), 0, 16) -- 6743
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(21,21),(13,13)), 0, 16) -- 6744
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(22,22),(14,14)), 0, 16) -- 6745
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(23,23),(15,15)), 0, 16) -- 6746
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(24,24),(16,16)), 0, 16) -- 6747
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(25,25),(17,17)), 0, 16) -- 6748
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(26,26),(18,18)), 0, 16) -- 6749
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 6750
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 6751
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 6752
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 6753
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 6754
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 6755
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 6756
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 6757
,( 5, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(18,18),(12,12)), 0, 16) -- 6758
,( 5, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(19,19),(13,13)), 0, 16) -- 6759
,( 5, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(20,20),(14,14)), 0, 16) -- 6760
,( 5, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(21,21),(15,15)), 0, 16) -- 6761
,( 5, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(22,22),(16,16)), 0, 16) -- 6762
,( 5, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(23,23),(17,17)), 0, 16) -- 6763
,( 5, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(24,24),(18,18)), 0, 16) -- 6764
,( 5, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(25,25),(19,19)), 0, 16) -- 6765
,( 5, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 6766
,( 5, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 6767
,( 5, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 6768
,( 5, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 6769
,( 5, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 6770
,( 5, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 6771
,( 5, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 6772
,( 5, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 6773
,( 5, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 6774
,( 5, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 6775
,( 5, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 6776
,( 5, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 6777
,( 5, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 6778
,( 5, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 6779
,( 5, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 6780
,( 5, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 6781
,( 5, E,0,0,((29,29),(99,99),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 6782
,( 5, E,0,0,((30,30),(99,99),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 6783
,( 5, E,0,0,((31,31),(99,99),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 6784
,( 5, E,0,0,((32,32),(99,99),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 6785
,( 5, E,0,0,((33,33),(99,99),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 6786
,( 5, E,0,0,((34,34),(99,99),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 6787
,( 5, E,0,0,((35,35),(99,99),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 6788
,( 5, E,0,0,((36,36),(99,99),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 6789
,( 5, E,0,0,((29,29),(99,99),( 0, 0),(17,17),(18,18),(10,10)), 0, 15) -- 6790
,( 5, E,0,0,((30,30),(99,99),( 1, 1),(18,18),(19,19),(11,11)), 0, 15) -- 6791
,( 5, E,0,0,((31,31),(99,99),( 2, 2),(19,19),(20,20),(12,12)), 0, 15) -- 6792
,( 5, E,0,0,((32,32),(99,99),( 3, 3),(20,20),(21,21),(13,13)), 0, 15) -- 6793
,( 5, E,0,0,((33,33),(99,99),( 4, 4),(21,21),(22,22),(14,14)), 0, 15) -- 6794
,( 5, E,0,0,((34,34),(99,99),( 5, 5),(22,22),(23,23),(15,15)), 0, 15) -- 6795
,( 5, E,0,0,((35,35),(99,99),( 6, 6),(23,23),(24,24),(16,16)), 0, 15) -- 6796
,( 5, E,0,0,((36,36),(99,99),( 7, 7),(24,24),(25,25),(17,17)), 0, 15) -- 6797
,( 5, E,0,0,((28,31),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 6798
,( 5, E,0,0,((30,33),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 6799
,( 5, E,0,0,((32,35),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 6800
,( 5, E,0,0,((34,37),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 6801
,( 5, E,0,0,((28,31),(23,23),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 6802
,( 5, E,0,0,((30,33),(25,25),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 6803
,( 5, E,0,0,((32,35),(27,27),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 6804
,( 5, E,0,0,((34,37),(29,29),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 6805
,( 5, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(20,21),(12,15)), 0, 13) -- 6806
,( 5, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(22,23),(14,17)), 0, 13) -- 6807
,( 5, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(24,25),(16,19)), 0, 13) -- 6808
,( 5, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(26,27),(18,21)), 0, 13) -- 6809
,( 5, E,0,0,((28,31),(23,23),( 0, 1),(18,19),(20,21),(10,13)), 0, 13) -- 6810
,( 5, E,0,0,((30,33),(25,25),( 2, 3),(20,21),(22,23),(12,15)), 0, 13) -- 6811
,( 5, E,0,0,((32,35),(27,27),( 4, 5),(22,23),(24,25),(14,17)), 0, 13) -- 6812
,( 5, E,0,0,((34,37),(29,29),( 6, 7),(24,25),(26,27),(16,19)), 0, 13) -- 6813
,( 5, E,0,0,((26,29),(22,22),( 0, 0),(16,17),(18,19),( 8,11)), 0, 13) -- 6814
,( 5, E,0,0,((28,31),(24,24),( 2, 2),(18,19),(20,21),(10,13)), 0, 13) -- 6815
,( 5, E,0,0,((30,33),(26,26),( 4, 4),(20,21),(22,23),(12,15)), 0, 13) -- 6816
,( 5, E,0,0,((32,35),(28,28),( 6, 6),(22,23),(24,25),(14,17)), 0, 13) -- 6817
,( 5, E,0,0,((26,29),(22,22),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 6818
,( 5, E,0,0,((28,31),(24,24),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 6819
,( 5, E,0,0,((30,33),(26,26),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 6820
,( 5, E,0,0,((32,35),(28,28),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 6821
,( 5, E,0,0,((26,27),(21,21),( 0, 0),(17,17),(19,19),(10,13)), 0, 12) -- 6822
,( 5, E,0,0,((28,29),(23,23),( 2, 2),(19,19),(21,21),(12,15)), 0, 12) -- 6823
,( 5, E,0,0,((30,31),(25,25),( 4, 4),(21,21),(23,23),(14,17)), 0, 12) -- 6824
,( 5, E,0,0,((32,33),(27,27),( 6, 6),(23,23),(25,25),(16,19)), 0, 12) -- 6825
,( 5, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(22,22),(14,17)), 0, 12) -- 6826
,( 5, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(24,24),(16,19)), 0, 12) -- 6827
,( 5, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(26,26),(18,21)), 0, 12) -- 6828
,( 5, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(28,28),(20,23)), 0, 12) -- 6829
,( 5, E,0,0,((26,29),(21,21),( 0, 1),(17,17),(20,20),(10,13)), 0, 12) -- 6830
,( 5, E,0,0,((28,31),(23,23),( 2, 3),(19,19),(22,22),(12,15)), 0, 12) -- 6831
,( 5, E,0,0,((30,33),(25,25),( 4, 5),(21,21),(24,24),(14,17)), 0, 12) -- 6832
,( 5, E,0,0,((32,35),(27,27),( 6, 7),(23,23),(26,26),(16,19)), 0, 12) -- 6833
,( 5, E,0,0,((24,27),(21,21),( 0, 1),(18,19),(20,21),(10,13)), 0, 11) -- 6834
,( 5, E,0,0,((26,29),(23,23),( 2, 3),(20,21),(22,23),(12,15)), 0, 11) -- 6835
,( 5, E,0,0,((28,31),(25,25),( 4, 5),(22,23),(24,25),(14,17)), 0, 11) -- 6836
,( 5, E,0,0,((30,33),(27,27),( 6, 7),(24,25),(26,27),(16,19)), 0, 11) -- 6837
,( 5, E,0,0,((24,25),(20,21),( 0, 0),(17,17),(20,21),(10,13)), 0, 11) -- 6838
,( 5, E,0,0,((26,27),(22,23),( 2, 2),(19,19),(22,23),(12,15)), 0, 11) -- 6839
,( 5, E,0,0,((28,29),(24,25),( 4, 4),(21,21),(24,25),(14,17)), 0, 11) -- 6840
,( 5, E,0,0,((30,31),(26,27),( 6, 6),(23,23),(26,27),(16,19)), 0, 11) -- 6841
,( 5, E,0,0,((24,27),(22,22),( 0, 1),(18,19),(22,23),(12,15)), 0, 11) -- 6842
,( 5, E,0,0,((26,29),(24,24),( 2, 3),(20,21),(24,25),(14,17)), 0, 11) -- 6843
,( 5, E,0,0,((28,31),(26,26),( 4, 5),(22,23),(26,27),(16,19)), 0, 11) -- 6844
,( 5, E,0,0,((30,33),(28,28),( 6, 7),(24,25),(28,29),(18,21)), 0, 11) -- 6845
,( 5, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 6846
,( 5, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 6847
,( 5, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 6848
,( 5, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 6849
,( 5, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 6850
,( 5, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 6851
,( 5, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 6852
,( 5, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 6853
,( 5, E,0,0,((26,29),(99,99),( 0, 1),(18,18),(19,19),( 8,11)), 0, 11) -- 6854
,( 5, E,0,0,((28,31),(99,99),( 2, 3),(20,20),(21,21),(10,13)), 0, 11) -- 6855
,( 5, E,0,0,((30,33),(99,99),( 4, 5),(22,22),(23,23),(12,15)), 0, 11) -- 6856
,( 5, E,0,0,((32,35),(99,99),( 6, 7),(24,24),(25,25),(14,17)), 0, 11) -- 6857
,( 5, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 6858
,( 5, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 6859
,( 5, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 6860
,( 5, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 6861
,( 5, E,0,0,((24,27),(21,21),( 0, 1),(16,17),(18,19),( 6, 9)), 0, 10) -- 6862
,( 5, E,0,0,((26,29),(23,23),( 2, 3),(18,19),(20,21),( 8,11)), 0, 10) -- 6863
,( 5, E,0,0,((28,31),(25,25),( 4, 5),(20,21),(22,23),(10,13)), 0, 10) -- 6864
,( 5, E,0,0,((30,33),(27,27),( 6, 7),(22,23),(24,25),(12,15)), 0, 10) -- 6865
,( 5, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(10,13)), 0, 10) -- 6866
,( 5, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(12,15)), 0, 10) -- 6867
,( 5, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(14,17)), 0, 10) -- 6868
,( 5, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(16,19)), 0, 10) -- 6869
,( 5, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 10) -- 6870
,( 5, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 10) -- 6871
,( 5, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 10) -- 6872
,( 5, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 10) -- 6873
,( 5, E,0,0,((24,27),(22,22),( 0, 1),(19,19),(22,22),( 8,11)), 0, 10) -- 6874
,( 5, E,0,0,((26,29),(24,24),( 2, 3),(21,21),(24,24),(10,13)), 0, 10) -- 6875
,( 5, E,0,0,((28,31),(26,26),( 4, 5),(23,23),(26,26),(12,15)), 0, 10) -- 6876
,( 5, E,0,0,((30,33),(28,28),( 6, 7),(25,25),(28,28),(14,17)), 0, 10) -- 6877
,( 5, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(18,19),( 4, 7)), 0, 10) -- 6878
,( 5, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(20,21),( 6, 9)), 0, 10) -- 6879
,( 5, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(22,23),( 8,11)), 0, 10) -- 6880
,( 5, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(24,25),(10,13)), 0, 10) -- 6881
,( 5, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,20),( 6, 9)), 0, 10) -- 6882
,( 5, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,22),( 8,11)), 0, 10) -- 6883
,( 5, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,24),(10,13)), 0, 10) -- 6884
,( 5, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,26),(12,15)), 0, 10) -- 6885
,( 5, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(18,19),( 2, 5)), 0, 10) -- 6886
,( 5, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(20,21),( 4, 7)), 0, 10) -- 6887
,( 5, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(22,23),( 6, 9)), 0, 10) -- 6888
,( 5, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(24,25),( 8,11)), 0, 10) -- 6889
,( 5, E,0,0,((22,23),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 10) -- 6890
,( 5, E,0,0,((24,25),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 10) -- 6891
,( 5, E,0,0,((26,27),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 10) -- 6892
,( 5, E,0,0,((28,29),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 10) -- 6893
,( 5, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 6894
,( 5, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 6895
,( 5, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 6896
,( 5, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 6897
,( 5, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 4, 7)), 0,  9) -- 6898
,( 5, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 6, 9)), 0,  9) -- 6899
,( 5, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 8,11)), 0,  9) -- 6900
,( 5, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),(10,13)), 0,  9) -- 6901
,( 5, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 6902
,( 5, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 6903
,( 5, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 6904
,( 5, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 6905
,( 5, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),( 6, 9)), 0,  9) -- 6906
,( 5, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),( 8,11)), 0,  9) -- 6907
,( 5, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(10,13)), 0,  9) -- 6908
,( 5, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(12,15)), 0,  9) -- 6909
,( 5, E,0,0,((20,23),(19,19),( 0, 1),(18,19),(20,21),( 8,11)), 0,  9) -- 6910
,( 5, E,0,0,((22,25),(21,21),( 2, 3),(20,21),(22,23),(10,13)), 0,  9) -- 6911
,( 5, E,0,0,((24,27),(23,23),( 4, 5),(22,23),(24,25),(12,15)), 0,  9) -- 6912
,( 5, E,0,0,((26,29),(25,25),( 6, 7),(24,25),(26,27),(14,17)), 0,  9) -- 6913
,( 5, E,0,0,((24,27),(21,21),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 6914
,( 5, E,0,0,((26,29),(23,23),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 6915
,( 5, E,0,0,((28,31),(25,25),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 6916
,( 5, E,0,0,((30,33),(27,27),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 6917
,( 5, E,0,0,((22,25),(20,21),( 1, 1),(20,21),(24,25),(14,17)), 0,  9) -- 6918
,( 5, E,0,0,((24,27),(22,23),( 3, 3),(22,23),(26,27),(16,19)), 0,  9) -- 6919
,( 5, E,0,0,((26,29),(24,25),( 5, 5),(24,25),(28,29),(18,21)), 0,  9) -- 6920
,( 5, E,0,0,((28,31),(26,27),( 7, 7),(26,27),(30,31),(20,23)), 0,  9) -- 6921
,( 5, E,0,0,((18,21),(18,19),( 0, 0),(18,19),(22,23),(10,13)), 0,  9) -- 6922
,( 5, E,0,0,((20,23),(20,21),( 2, 2),(20,21),(24,25),(12,15)), 0,  9) -- 6923
,( 5, E,0,0,((22,25),(22,23),( 4, 4),(22,23),(26,27),(14,17)), 0,  9) -- 6924
,( 5, E,0,0,((24,27),(24,25),( 6, 6),(24,25),(28,29),(16,19)), 0,  9) -- 6925
,( 5, E,0,0,((20,23),(20,21),( 0, 1),(20,20),(22,23),(14,15)), 0,  9) -- 6926
,( 5, E,0,0,((22,25),(22,23),( 2, 3),(22,22),(24,25),(16,17)), 0,  9) -- 6927
,( 5, E,0,0,((24,27),(24,25),( 4, 5),(24,24),(26,27),(18,19)), 0,  9) -- 6928
,( 5, E,0,0,((26,29),(26,27),( 6, 7),(26,26),(28,29),(20,21)), 0,  9) -- 6929
,( 5, E,0,0,((20,23),(20,21),( 0, 0),(18,18),(20,21),(10,11)), 0,  9) -- 6930
,( 5, E,0,0,((22,25),(22,23),( 2, 2),(20,20),(22,23),(12,13)), 0,  9) -- 6931
,( 5, E,0,0,((24,27),(24,25),( 4, 4),(22,22),(24,25),(14,15)), 0,  9) -- 6932
,( 5, E,0,0,((26,29),(26,27),( 6, 6),(24,24),(26,27),(16,17)), 0,  9) -- 6933
,( 5, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),( 6, 9)), 0,  9) -- 6934
,( 5, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),( 8,11)), 0,  9) -- 6935
,( 5, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(10,13)), 0,  9) -- 6936
,( 5, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(12,15)), 0,  9) -- 6937
,( 5, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(24,25),(10,13)), 0,  9) -- 6938
,( 5, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(26,27),(12,15)), 0,  9) -- 6939
,( 5, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(28,29),(14,17)), 0,  9) -- 6940
,( 5, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(30,31),(16,19)), 0,  9) -- 6941
,( 5, E,0,0,((23,23),(20,21),( 0, 0),(18,18),(20,21),( 2, 5)), 0,  9) -- 6942
,( 5, E,0,0,((25,25),(22,23),( 2, 2),(20,20),(22,23),( 4, 7)), 0,  9) -- 6943
,( 5, E,0,0,((27,27),(24,25),( 4, 4),(22,22),(24,25),( 6, 9)), 0,  9) -- 6944
,( 5, E,0,0,((29,29),(26,27),( 6, 6),(24,24),(26,27),( 8,11)), 0,  9) -- 6945
,( 5, E,0,0,((24,25),(22,22),( 1, 1),(18,19),(20,21),( 8,11)), 0,  9) -- 6946
,( 5, E,0,0,((26,27),(24,24),( 3, 3),(20,21),(22,23),(10,13)), 0,  9) -- 6947
,( 5, E,0,0,((28,29),(26,26),( 5, 5),(22,23),(24,25),(12,15)), 0,  9) -- 6948
,( 5, E,0,0,((30,31),(28,28),( 7, 7),(24,25),(26,27),(14,17)), 0,  9) -- 6949
,( 5, E,0,0,((24,27),(21,21),( 1, 1),(20,20),(22,23),(12,15)), 0,  9) -- 6950
,( 5, E,0,0,((26,29),(23,23),( 3, 3),(22,22),(24,25),(14,17)), 0,  9) -- 6951
,( 5, E,0,0,((28,31),(25,25),( 5, 5),(24,24),(26,27),(16,19)), 0,  9) -- 6952
,( 5, E,0,0,((30,33),(27,27),( 7, 7),(26,26),(28,29),(18,21)), 0,  9) -- 6953
,( 5, E,0,0,((20,23),(20,21),( 1, 1),(20,21),(24,24),( 6, 9)), 0,  9) -- 6954
,( 5, E,0,0,((22,25),(22,23),( 3, 3),(22,23),(26,26),( 8,11)), 0,  9) -- 6955
,( 5, E,0,0,((24,27),(24,25),( 5, 5),(24,25),(28,28),(10,13)), 0,  9) -- 6956
,( 5, E,0,0,((26,29),(26,27),( 7, 7),(26,27),(30,30),(12,15)), 0,  9) -- 6957
,( 5, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(18,19),( 1, 1)), 0,  9) -- 6958
,( 5, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(20,21),( 3, 3)), 0,  9) -- 6959
,( 5, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(22,23),( 5, 5)), 0,  9) -- 6960
,( 5, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(24,25),( 7, 7)), 0,  9) -- 6961
,( 5, E,0,0,((20,23),(19,19),( 0, 1),(19,19),(22,23),( 4, 7)), 0,  9) -- 6962
,( 5, E,0,0,((22,25),(21,21),( 2, 3),(21,21),(24,25),( 6, 9)), 0,  9) -- 6963
,( 5, E,0,0,((24,27),(23,23),( 4, 5),(23,23),(26,27),( 8,11)), 0,  9) -- 6964
,( 5, E,0,0,((26,29),(25,25),( 6, 7),(25,25),(28,29),(10,13)), 0,  9) -- 6965
,( 5, E,0,0,((24,27),(22,22),( 0, 1),(18,18),(19,19),( 0, 3)), 0,  9) -- 6966
,( 5, E,0,0,((26,29),(24,24),( 2, 3),(20,20),(21,21),( 2, 5)), 0,  9) -- 6967
,( 5, E,0,0,((28,31),(26,26),( 4, 5),(22,22),(23,23),( 4, 7)), 0,  9) -- 6968
,( 5, E,0,0,((30,33),(28,28),( 6, 7),(24,24),(25,25),( 6, 9)), 0,  9) -- 6969
,( 5, E,0,0,((22,25),(99,99),( 1, 1),(20,20),(20,21),( 8, 8)), 0,  9) -- 6970
,( 5, E,0,0,((24,27),(99,99),( 3, 3),(22,22),(22,23),(10,10)), 0,  9) -- 6971
,( 5, E,0,0,((26,29),(99,99),( 5, 5),(24,24),(24,25),(12,12)), 0,  9) -- 6972
,( 5, E,0,0,((28,31),(99,99),( 7, 7),(26,26),(26,27),(14,14)), 0,  9) -- 6973
,( 5, E,0,0,((24,27),(99,99),( 0, 1),(16,17),(16,17),(99,99)), 0,  9) -- 6974
,( 5, E,0,0,((26,29),(99,99),( 2, 3),(18,19),(18,19),(99,99)), 0,  9) -- 6975
,( 5, E,0,0,((28,31),(99,99),( 4, 5),(20,21),(20,21),(99,99)), 0,  9) -- 6976
,( 5, E,0,0,((30,33),(99,99),( 6, 7),(22,23),(22,23),(99,99)), 0,  9) -- 6977
,( 5, E,0,0,((18,21),(18,21),( 0, 1),(18,21),(18,21),(99,99)), 0,  8) -- 6978
,( 5, E,0,0,((20,23),(20,23),( 2, 3),(20,23),(20,23),(99,99)), 0,  8) -- 6979
,( 5, E,0,0,((22,25),(22,25),( 4, 5),(22,25),(22,25),(99,99)), 0,  8) -- 6980
,( 5, E,0,0,((24,27),(24,27),( 6, 7),(24,27),(24,27),(99,99)), 0,  8) -- 6981
,( 5, E,0,0,((18,21),(18,21),( 0, 1),(18,21),(22,25),(99,99)), 0,  8) -- 6982
,( 5, E,0,0,((20,23),(20,23),( 2, 3),(20,23),(24,27),(99,99)), 0,  8) -- 6983
,( 5, E,0,0,((22,25),(22,25),( 4, 5),(22,25),(26,29),(99,99)), 0,  8) -- 6984
,( 5, E,0,0,((24,27),(24,27),( 6, 7),(24,27),(28,31),(99,99)), 0,  8) -- 6985
,( 5, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 6986
,( 5, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 6987
,( 5, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 6988
,( 5, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 6989
,( 5, E,0,0,((14,17),(16,19),( 0, 1),(18,21),(20,23),(99,99)), 0,  7) -- 6990
,( 5, E,0,0,((16,19),(18,21),( 2, 3),(20,23),(22,25),(99,99)), 0,  7) -- 6991
,( 5, E,0,0,((18,21),(20,23),( 4, 5),(22,25),(24,27),(99,99)), 0,  7) -- 6992
,( 5, E,0,0,((20,23),(22,25),( 6, 7),(24,27),(26,29),(99,99)), 0,  7) -- 6993
,( 5, E,0,1,((16,19),(16,19),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 6994
,( 5, E,0,1,((18,21),(18,21),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 6995
,( 5, E,0,1,((20,23),(20,23),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 6996
,( 5, E,0,1,((22,25),(22,25),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 6997
,( 5, E,0,1,((12,15),(16,19),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 6998
,( 5, E,0,1,((14,17),(18,21),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 6999
,( 5, E,0,1,((16,19),(20,23),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 7000
,( 5, E,0,1,((18,21),(22,25),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 7001
,( 5, E,0,1,((16,19),(18,21),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 7002
,( 5, E,0,1,((18,21),(20,23),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 7003
,( 5, E,0,1,((20,23),(22,25),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 7004
,( 5, E,0,1,((22,25),(24,27),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 7005
,( 5, E,0,1,((20,23),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 7006
,( 5, E,0,1,((22,25),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 7007
,( 5, E,0,1,((24,27),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 7008
,( 5, E,0,1,((26,29),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 7009
,( 5, E,0,1,((20,23),(99,99),( 0, 1),(20,21),(99,99),(99,99)), 0,  7) -- 7010
,( 5, E,0,1,((22,25),(99,99),( 2, 3),(22,23),(99,99),(99,99)), 0,  7) -- 7011
,( 5, E,0,1,((24,27),(99,99),( 4, 5),(24,25),(99,99),(99,99)), 0,  7) -- 7012
,( 5, E,0,1,((26,29),(99,99),( 6, 7),(26,27),(99,99),(99,99)), 0,  7) -- 7013
,( 5, E,0,1,((24,27),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 7014
,( 5, E,0,1,((26,29),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 7015
,( 5, E,0,1,((28,31),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 7016
,( 5, E,0,1,((30,33),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 7017
,( 5, E,0,1,((20,23),(20,23),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 7018
,( 5, E,0,1,((22,25),(22,25),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 7019
,( 5, E,0,1,((24,27),(24,27),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 7020
,( 5, E,0,1,((26,29),(26,29),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 7021
,( 5, E,0,1,((24,27),(22,22),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 7022
,( 5, E,0,1,((26,29),(24,24),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 7023
,( 5, E,0,1,((28,31),(26,26),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 7024
,( 5, E,0,1,((30,33),(28,28),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 7025
,( 5, E,0,1,(( 8,11),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  6) -- 7026
,( 5, E,0,1,((10,13),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  6) -- 7027
,( 5, E,0,1,((12,15),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  6) -- 7028
,( 5, E,0,1,((14,17),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  6) -- 7029
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 7030
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 7031
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 7032
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 7033
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 7034
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 7035
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 7036
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 7037
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 31) -- 7038
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 31) -- 7039
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 31) -- 7040
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 31) -- 7041
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 31) -- 7042
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 31) -- 7043
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 31) -- 7044
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 31) -- 7045
,( 6, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 30) -- 7046
,( 6, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 30) -- 7047
,( 6, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 30) -- 7048
,( 6, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 30) -- 7049
,( 6, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 30) -- 7050
,( 6, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 30) -- 7051
,( 6, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 30) -- 7052
,( 6, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 30) -- 7053
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 30) -- 7054
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 30) -- 7055
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 30) -- 7056
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 30) -- 7057
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 30) -- 7058
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 30) -- 7059
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 30) -- 7060
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 30) -- 7061
,( 6, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 30) -- 7062
,( 6, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 30) -- 7063
,( 6, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 30) -- 7064
,( 6, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 30) -- 7065
,( 6, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 30) -- 7066
,( 6, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 30) -- 7067
,( 6, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 30) -- 7068
,( 6, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 30) -- 7069
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 28) -- 7070
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 28) -- 7071
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 28) -- 7072
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 28) -- 7073
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 28) -- 7074
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 28) -- 7075
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 28) -- 7076
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 28) -- 7077
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 27) -- 7078
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 27) -- 7079
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 27) -- 7080
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 27) -- 7081
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 27) -- 7082
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 27) -- 7083
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 27) -- 7084
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 27) -- 7085
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 26) -- 7086
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 26) -- 7087
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 26) -- 7088
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 26) -- 7089
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 26) -- 7090
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 26) -- 7091
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 26) -- 7092
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 26) -- 7093
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 25) -- 7094
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 25) -- 7095
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 25) -- 7096
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 25) -- 7097
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 25) -- 7098
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 25) -- 7099
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 25) -- 7100
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 25) -- 7101
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 25) -- 7102
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 25) -- 7103
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),(10,10)), 1, 25) -- 7104
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(11,11)), 1, 25) -- 7105
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(12,12)), 1, 25) -- 7106
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(13,13)), 1, 25) -- 7107
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(14,14)), 1, 25) -- 7108
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(15,15)), 1, 25) -- 7109
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 24) -- 7110
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 24) -- 7111
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 24) -- 7112
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 24) -- 7113
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 24) -- 7114
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 24) -- 7115
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 24) -- 7116
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 24) -- 7117
,( 6, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 24) -- 7118
,( 6, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 24) -- 7119
,( 6, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 24) -- 7120
,( 6, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 24) -- 7121
,( 6, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 24) -- 7122
,( 6, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 24) -- 7123
,( 6, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 24) -- 7124
,( 6, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 24) -- 7125
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 7126
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 7127
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 7128
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 7129
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 7130
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 7131
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 7132
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 7133
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 22) -- 7134
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 22) -- 7135
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 22) -- 7136
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 22) -- 7137
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 22) -- 7138
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 22) -- 7139
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 22) -- 7140
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 22) -- 7141
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 21) -- 7142
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 21) -- 7143
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 21) -- 7144
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 21) -- 7145
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 21) -- 7146
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 21) -- 7147
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 21) -- 7148
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 21) -- 7149
,( 6, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 21) -- 7150
,( 6, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 21) -- 7151
,( 6, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 21) -- 7152
,( 6, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 21) -- 7153
,( 6, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 21) -- 7154
,( 6, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 21) -- 7155
,( 6, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 21) -- 7156
,( 6, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 21) -- 7157
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 20) -- 7158
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 20) -- 7159
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 20) -- 7160
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 20) -- 7161
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 20) -- 7162
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 20) -- 7163
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 20) -- 7164
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 20) -- 7165
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 20) -- 7166
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 20) -- 7167
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 20) -- 7168
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 20) -- 7169
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 20) -- 7170
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 20) -- 7171
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 20) -- 7172
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 20) -- 7173
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 8, 8)), 1, 20) -- 7174
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 9, 9)), 1, 20) -- 7175
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),(10,10)), 1, 20) -- 7176
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(11,11)), 1, 20) -- 7177
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(12,12)), 1, 20) -- 7178
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(13,13)), 1, 20) -- 7179
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(14,14)), 1, 20) -- 7180
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(15,15)), 1, 20) -- 7181
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 19) -- 7182
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 19) -- 7183
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 19) -- 7184
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(19,19),(18,18),(10,10)), 1, 19) -- 7185
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(20,20),(19,19),(11,11)), 1, 19) -- 7186
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(21,21),(20,20),(12,12)), 1, 19) -- 7187
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(22,22),(21,21),(13,13)), 1, 19) -- 7188
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(23,23),(22,22),(14,14)), 1, 19) -- 7189
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 7190
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 7191
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 7192
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 7193
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 7194
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 7195
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 7196
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 7197
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 19) -- 7198
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 19) -- 7199
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 19) -- 7200
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 19) -- 7201
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 19) -- 7202
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 19) -- 7203
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 19) -- 7204
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 19) -- 7205
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(16,16),(15,15),( 6, 6)), 1, 19) -- 7206
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(17,17),(16,16),( 7, 7)), 1, 19) -- 7207
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(18,18),(17,17),( 8, 8)), 1, 19) -- 7208
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(19,19),(18,18),( 9, 9)), 1, 19) -- 7209
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(20,20),(19,19),(10,10)), 1, 19) -- 7210
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(21,21),(20,20),(11,11)), 1, 19) -- 7211
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(22,22),(21,21),(12,12)), 1, 19) -- 7212
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(23,23),(22,22),(13,13)), 1, 19) -- 7213
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 7214
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 7215
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 7216
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 7217
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 7218
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 7219
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 7220
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 7221
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 7222
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 7223
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 7224
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 7225
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 7226
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 7227
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 7228
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 7229
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 7230
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 7231
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 7232
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 7233
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 7234
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 7235
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 7236
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 7237
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 7238
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 7239
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 7240
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 7241
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 7242
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 7243
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 7244
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 7245
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 7246
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 7247
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 7248
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 7249
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 7250
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 7251
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 7252
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 7253
,( 6, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 18) -- 7254
,( 6, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 18) -- 7255
,( 6, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 18) -- 7256
,( 6, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 18) -- 7257
,( 6, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 18) -- 7258
,( 6, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 18) -- 7259
,( 6, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 18) -- 7260
,( 6, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 18) -- 7261
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 7262
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 7263
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 7264
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 7265
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 7266
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 7267
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 7268
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 7269
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 7270
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 7271
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 7272
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 7273
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 7274
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 7275
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 7276
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 7277
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 7278
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 7279
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 7280
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 7281
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 7282
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 7283
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 7284
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 7285
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 17) -- 7286
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 17) -- 7287
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 17) -- 7288
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 17) -- 7289
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 17) -- 7290
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 17) -- 7291
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 17) -- 7292
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 17) -- 7293
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 7294
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 7295
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 7296
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 7297
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 7298
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 7299
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 7300
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 7301
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 16) -- 7302
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 16) -- 7303
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 16) -- 7304
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 16) -- 7305
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 16) -- 7306
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 16) -- 7307
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 16) -- 7308
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 16) -- 7309
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 16) -- 7310
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 16) -- 7311
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 16) -- 7312
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 16) -- 7313
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 16) -- 7314
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 16) -- 7315
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 16) -- 7316
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 16) -- 7317
,( 6, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 16) -- 7318
,( 6, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 16) -- 7319
,( 6, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 16) -- 7320
,( 6, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 16) -- 7321
,( 6, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 16) -- 7322
,( 6, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 16) -- 7323
,( 6, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 16) -- 7324
,( 6, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 16) -- 7325
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(13,13),( 4, 4)), 1, 16) -- 7326
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(14,14),( 5, 5)), 1, 16) -- 7327
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(15,15),( 6, 6)), 1, 16) -- 7328
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(16,16),( 7, 7)), 1, 16) -- 7329
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(17,17),( 8, 8)), 1, 16) -- 7330
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(18,18),( 9, 9)), 1, 16) -- 7331
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(19,19),(10,10)), 1, 16) -- 7332
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(20,20),(11,11)), 1, 16) -- 7333
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 16) -- 7334
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 16) -- 7335
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 16) -- 7336
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 16) -- 7337
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 16) -- 7338
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 16) -- 7339
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 16) -- 7340
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 16) -- 7341
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 16) -- 7342
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 16) -- 7343
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 16) -- 7344
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),(10,10)), 1, 16) -- 7345
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(11,11)), 1, 16) -- 7346
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(12,12)), 1, 16) -- 7347
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(13,13)), 1, 16) -- 7348
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(14,14)), 1, 16) -- 7349
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 7350
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 7351
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 7352
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 7353
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 7354
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 7355
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 7356
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 7357
,( 6, E,0,0,((36,36),(99,99),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 16) -- 7358
,( 6, E,0,0,((37,37),(99,99),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 16) -- 7359
,( 6, E,0,0,((38,38),(99,99),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 16) -- 7360
,( 6, E,0,0,((39,39),(99,99),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 16) -- 7361
,( 6, E,0,0,((40,40),(99,99),( 4, 4),(19,19),(19,19),(10,10)), 1, 16) -- 7362
,( 6, E,0,0,((41,41),(99,99),( 5, 5),(20,20),(20,20),(11,11)), 1, 16) -- 7363
,( 6, E,0,0,((42,42),(99,99),( 6, 6),(21,21),(21,21),(12,12)), 1, 16) -- 7364
,( 6, E,0,0,((43,43),(99,99),( 7, 7),(22,22),(22,22),(13,13)), 1, 16) -- 7365
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 7366
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 7367
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 7368
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 7369
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 7370
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 7371
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 7372
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 7373
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 15) -- 7374
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 15) -- 7375
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 15) -- 7376
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 15) -- 7377
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 15) -- 7378
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(18,18),(10,10)), 1, 15) -- 7379
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(19,19),(11,11)), 1, 15) -- 7380
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(20,20),(12,12)), 1, 15) -- 7381
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 15) -- 7382
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 15) -- 7383
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 15) -- 7384
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),(10,10)), 1, 15) -- 7385
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),(11,11)), 1, 15) -- 7386
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(12,12)), 1, 15) -- 7387
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(13,13)), 1, 15) -- 7388
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(14,14)), 1, 15) -- 7389
,( 6, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 7390
,( 6, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 7391
,( 6, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 7392
,( 6, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 7393
,( 6, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 7394
,( 6, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 7395
,( 6, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 7396
,( 6, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 7397
,( 6, E,0,0,((36,36),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 7398
,( 6, E,0,0,((37,37),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 7399
,( 6, E,0,0,((38,38),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 7400
,( 6, E,0,0,((39,39),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 7401
,( 6, E,0,0,((40,40),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 7402
,( 6, E,0,0,((41,41),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 7403
,( 6, E,0,0,((42,42),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 7404
,( 6, E,0,0,((43,43),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 7405
,( 6, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 7406
,( 6, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 7407
,( 6, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 7408
,( 6, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 7409
,( 6, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 7410
,( 6, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 7411
,( 6, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 7412
,( 6, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 7413
,( 6, E,0,0,((36,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 7414
,( 6, E,0,0,((38,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 7415
,( 6, E,0,0,((40,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 7416
,( 6, E,0,0,((42,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 7417
,( 6, E,0,0,((38,41),(28,29),( 1, 1),(15,15),(14,14),( 4, 7)), 1, 13) -- 7418
,( 6, E,0,0,((40,43),(30,31),( 3, 3),(17,17),(16,16),( 6, 9)), 1, 13) -- 7419
,( 6, E,0,0,((42,45),(32,33),( 5, 5),(19,19),(18,18),( 8,11)), 1, 13) -- 7420
,( 6, E,0,0,((44,47),(34,35),( 7, 7),(21,21),(20,20),(10,13)), 1, 13) -- 7421
,( 6, E,0,0,((36,39),(28,29),( 0, 1),(14,15),(12,13),( 4, 7)), 1, 13) -- 7422
,( 6, E,0,0,((38,41),(30,31),( 2, 3),(16,17),(14,15),( 6, 9)), 1, 13) -- 7423
,( 6, E,0,0,((40,43),(32,33),( 4, 5),(18,19),(16,17),( 8,11)), 1, 13) -- 7424
,( 6, E,0,0,((42,45),(34,35),( 6, 7),(20,21),(18,19),(10,13)), 1, 13) -- 7425
,( 6, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 7426
,( 6, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 7427
,( 6, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 7428
,( 6, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 7429
,( 6, E,0,0,((36,39),(26,27),( 0, 0),(14,15),(12,13),( 6, 9)), 1, 12) -- 7430
,( 6, E,0,0,((38,41),(28,29),( 2, 2),(16,17),(14,15),( 8,11)), 1, 12) -- 7431
,( 6, E,0,0,((40,43),(30,31),( 4, 4),(18,19),(16,17),(10,13)), 1, 12) -- 7432
,( 6, E,0,0,((42,45),(32,33),( 6, 6),(20,21),(18,19),(12,15)), 1, 12) -- 7433
,( 6, E,0,0,((38,41),(28,29),( 1, 1),(16,16),(14,15),( 6, 9)), 1, 12) -- 7434
,( 6, E,0,0,((40,43),(30,31),( 3, 3),(18,18),(16,17),( 8,11)), 1, 12) -- 7435
,( 6, E,0,0,((42,45),(32,33),( 5, 5),(20,20),(18,19),(10,13)), 1, 12) -- 7436
,( 6, E,0,0,((44,47),(34,35),( 7, 7),(22,22),(20,21),(12,15)), 1, 12) -- 7437
,( 6, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 12) -- 7438
,( 6, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 12) -- 7439
,( 6, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 12) -- 7440
,( 6, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 12) -- 7441
,( 6, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 7442
,( 6, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 7443
,( 6, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 7444
,( 6, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 7445
,( 6, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 11) -- 7446
,( 6, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 11) -- 7447
,( 6, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 11) -- 7448
,( 6, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 11) -- 7449
,( 6, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(10,11),( 0, 3)), 1, 11) -- 7450
,( 6, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(12,13),( 2, 5)), 1, 11) -- 7451
,( 6, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(14,15),( 4, 7)), 1, 11) -- 7452
,( 6, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(16,17),( 6, 9)), 1, 11) -- 7453
,( 6, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 8,11)), 1, 11) -- 7454
,( 6, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(10,13)), 1, 11) -- 7455
,( 6, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(12,15)), 1, 11) -- 7456
,( 6, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(14,17)), 1, 11) -- 7457
,( 6, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 7458
,( 6, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 7459
,( 6, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 7460
,( 6, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 7461
,( 6, E,0,0,((38,41),(27,27),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 11) -- 7462
,( 6, E,0,0,((40,43),(29,29),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 11) -- 7463
,( 6, E,0,0,((42,45),(31,31),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 11) -- 7464
,( 6, E,0,0,((44,47),(33,33),( 6, 6),(19,19),(18,18),( 8,11)), 1, 11) -- 7465
,( 6, E,0,0,((38,41),(28,28),( 0, 0),(13,13),(10,11),( 4, 5)), 1, 11) -- 7466
,( 6, E,0,0,((40,43),(30,30),( 2, 2),(15,15),(12,13),( 6, 7)), 1, 11) -- 7467
,( 6, E,0,0,((42,45),(32,32),( 4, 4),(17,17),(14,15),( 8, 9)), 1, 11) -- 7468
,( 6, E,0,0,((44,47),(34,34),( 6, 6),(19,19),(16,17),(10,11)), 1, 11) -- 7469
,( 6, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(10,11),( 2, 5)), 1, 10) -- 7470
,( 6, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(12,13),( 4, 7)), 1, 10) -- 7471
,( 6, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(14,15),( 6, 9)), 1, 10) -- 7472
,( 6, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(16,17),( 8,11)), 1, 10) -- 7473
,( 6, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 7474
,( 6, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 7475
,( 6, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(10,13)), 1, 10) -- 7476
,( 6, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(12,15)), 1, 10) -- 7477
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(10,11),( 2, 5)), 1, 10) -- 7478
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(12,13),( 4, 7)), 1, 10) -- 7479
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(14,15),( 6, 9)), 1, 10) -- 7480
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(16,17),( 8,11)), 1, 10) -- 7481
,( 6, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),( 6, 9)), 1, 10) -- 7482
,( 6, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),( 8,11)), 1, 10) -- 7483
,( 6, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(10,13)), 1, 10) -- 7484
,( 6, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(12,15)), 1, 10) -- 7485
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1, 10) -- 7486
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1, 10) -- 7487
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 8,11)), 1, 10) -- 7488
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(10,13)), 1, 10) -- 7489
,( 6, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 7490
,( 6, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 7491
,( 6, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 7492
,( 6, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 7493
,( 6, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1, 10) -- 7494
,( 6, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 8,11)), 1, 10) -- 7495
,( 6, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(10,13)), 1, 10) -- 7496
,( 6, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(12,15)), 1, 10) -- 7497
,( 6, E,0,0,((42,43),(30,30),( 1, 1),(14,15),(14,14),( 6, 9)), 1, 10) -- 7498
,( 6, E,0,0,((44,45),(32,32),( 3, 3),(16,17),(16,16),( 8,11)), 1, 10) -- 7499
,( 6, E,0,0,((46,47),(34,34),( 5, 5),(18,19),(18,18),(10,13)), 1, 10) -- 7500
,( 6, E,0,0,((48,49),(36,36),( 7, 7),(20,21),(20,20),(12,15)), 1, 10) -- 7501
,( 6, E,0,0,((40,43),(30,30),( 0, 1),(14,15),(12,13),(10,13)), 1, 10) -- 7502
,( 6, E,0,0,((42,45),(32,32),( 2, 3),(16,17),(14,15),(12,15)), 1, 10) -- 7503
,( 6, E,0,0,((44,47),(34,34),( 4, 5),(18,19),(16,17),(14,17)), 1, 10) -- 7504
,( 6, E,0,0,((46,49),(36,36),( 6, 7),(20,21),(18,19),(16,19)), 1, 10) -- 7505
,( 6, E,0,0,((40,43),(28,29),( 0, 0),(12,13),( 9, 9),( 0, 1)), 1, 10) -- 7506
,( 6, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(11,11),( 2, 3)), 1, 10) -- 7507
,( 6, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(13,13),( 4, 5)), 1, 10) -- 7508
,( 6, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(15,15),( 6, 7)), 1, 10) -- 7509
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1, 10) -- 7510
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1, 10) -- 7511
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1, 10) -- 7512
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1, 10) -- 7513
,( 6, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,12),( 4, 5)), 1, 10) -- 7514
,( 6, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,14),( 6, 7)), 1, 10) -- 7515
,( 6, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,16),( 8, 9)), 1, 10) -- 7516
,( 6, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,18),(10,11)), 1, 10) -- 7517
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 8,11)), 1,  9) -- 7518
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),(10,13)), 1,  9) -- 7519
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(12,15)), 1,  9) -- 7520
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(14,17)), 1,  9) -- 7521
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 7522
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 7523
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 7524
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 7525
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 8,11)), 1,  9) -- 7526
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(10,13)), 1,  9) -- 7527
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(12,15)), 1,  9) -- 7528
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(14,17)), 1,  9) -- 7529
,( 6, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(12,13),(10,13)), 1,  9) -- 7530
,( 6, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(14,15),(12,15)), 1,  9) -- 7531
,( 6, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(16,17),(14,17)), 1,  9) -- 7532
,( 6, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(18,19),(16,19)), 1,  9) -- 7533
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),(10,13)), 1,  9) -- 7534
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(12,15)), 1,  9) -- 7535
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(14,17)), 1,  9) -- 7536
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(16,19)), 1,  9) -- 7537
,( 6, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(14,15),(12,15)), 1,  9) -- 7538
,( 6, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(16,17),(14,17)), 1,  9) -- 7539
,( 6, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(18,19),(16,19)), 1,  9) -- 7540
,( 6, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(20,21),(18,21)), 1,  9) -- 7541
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 0, 3)), 1,  9) -- 7542
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 2, 5)), 1,  9) -- 7543
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 4, 7)), 1,  9) -- 7544
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 6, 9)), 1,  9) -- 7545
,( 6, E,0,0,((46,49),(32,33),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 7546
,( 6, E,0,0,((48,51),(34,35),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 7547
,( 6, E,0,0,((50,53),(36,37),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 7548
,( 6, E,0,0,((52,55),(38,39),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 7549
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(11,11),( 6, 9)), 1,  9) -- 7550
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(13,13),( 8,11)), 1,  9) -- 7551
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(15,15),(10,13)), 1,  9) -- 7552
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(17,17),(12,15)), 1,  9) -- 7553
,( 6, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(12,13),(10,13)), 1,  9) -- 7554
,( 6, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(14,15),(12,15)), 1,  9) -- 7555
,( 6, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(16,17),(14,17)), 1,  9) -- 7556
,( 6, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(18,19),(16,19)), 1,  9) -- 7557
,( 6, E,0,0,((44,47),(30,31),( 0, 1),(12,13),( 8, 9),( 4, 7)), 1,  9) -- 7558
,( 6, E,0,0,((46,49),(32,33),( 2, 3),(14,15),(10,11),( 6, 9)), 1,  9) -- 7559
,( 6, E,0,0,((48,51),(34,35),( 4, 5),(16,17),(12,13),( 8,11)), 1,  9) -- 7560
,( 6, E,0,0,((50,53),(36,37),( 6, 7),(18,19),(14,15),(10,13)), 1,  9) -- 7561
,( 6, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(12,12),( 4, 7)), 1,  9) -- 7562
,( 6, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(14,14),( 6, 9)), 1,  9) -- 7563
,( 6, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(16,16),( 8,11)), 1,  9) -- 7564
,( 6, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(18,18),(10,13)), 1,  9) -- 7565
,( 6, E,0,0,((44,47),(32,32),( 1, 1),(14,14),(10,11),( 2, 5)), 1,  9) -- 7566
,( 6, E,0,0,((46,49),(34,34),( 3, 3),(16,16),(12,13),( 4, 7)), 1,  9) -- 7567
,( 6, E,0,0,((48,51),(36,36),( 5, 5),(18,18),(14,15),( 6, 9)), 1,  9) -- 7568
,( 6, E,0,0,((50,53),(38,38),( 7, 7),(20,20),(16,17),( 8,11)), 1,  9) -- 7569
,( 6, E,0,0,((44,47),(32,32),( 1, 1),(14,14),(12,13),( 8, 9)), 1,  9) -- 7570
,( 6, E,0,0,((46,49),(34,34),( 3, 3),(16,16),(14,15),(10,11)), 1,  9) -- 7571
,( 6, E,0,0,((48,51),(36,36),( 5, 5),(18,18),(16,17),(12,13)), 1,  9) -- 7572
,( 6, E,0,0,((50,53),(38,38),( 7, 7),(20,20),(18,19),(14,15)), 1,  9) -- 7573
,( 6, E,0,0,((44,47),(30,31),( 0, 1),(13,13),(12,12),( 6, 9)), 1,  9) -- 7574
,( 6, E,0,0,((46,49),(32,33),( 2, 3),(15,15),(14,14),( 8,11)), 1,  9) -- 7575
,( 6, E,0,0,((48,51),(34,35),( 4, 5),(17,17),(16,16),(10,13)), 1,  9) -- 7576
,( 6, E,0,0,((50,53),(36,37),( 6, 7),(19,19),(18,18),(12,15)), 1,  9) -- 7577
,( 6, E,0,0,((42,45),(30,30),( 1, 1),(14,15),(14,15),(14,17)), 1,  9) -- 7578
,( 6, E,0,0,((44,47),(32,32),( 3, 3),(16,17),(16,17),(16,19)), 1,  9) -- 7579
,( 6, E,0,0,((46,49),(34,34),( 5, 5),(18,19),(18,19),(18,21)), 1,  9) -- 7580
,( 6, E,0,0,((48,51),(36,36),( 7, 7),(20,21),(20,21),(20,23)), 1,  9) -- 7581
,( 6, E,0,0,((44,47),(31,31),( 0, 1),(12,13),(10,11),(10,13)), 1,  9) -- 7582
,( 6, E,0,0,((46,49),(33,33),( 2, 3),(14,15),(12,13),(12,15)), 1,  9) -- 7583
,( 6, E,0,0,((48,51),(35,35),( 4, 5),(16,17),(14,15),(14,17)), 1,  9) -- 7584
,( 6, E,0,0,((50,53),(37,37),( 6, 7),(18,19),(16,17),(16,19)), 1,  9) -- 7585
,( 6, E,0,0,((42,43),(28,29),( 0, 0),(13,13),(14,15),(14,17)), 1,  9) -- 7586
,( 6, E,0,0,((44,45),(30,31),( 2, 2),(15,15),(16,17),(16,19)), 1,  9) -- 7587
,( 6, E,0,0,((46,47),(32,33),( 4, 4),(17,17),(18,19),(18,21)), 1,  9) -- 7588
,( 6, E,0,0,((48,49),(34,35),( 6, 6),(19,19),(20,21),(20,23)), 1,  9) -- 7589
,( 6, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(12,15),( 8,11)), 1,  8) -- 7590
,( 6, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(14,17),(10,13)), 1,  8) -- 7591
,( 6, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(16,19),(12,15)), 1,  8) -- 7592
,( 6, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(18,21),(14,17)), 1,  8) -- 7593
,( 6, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(12,15)), 1,  8) -- 7594
,( 6, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(14,17)), 1,  8) -- 7595
,( 6, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(16,19)), 1,  8) -- 7596
,( 6, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(18,21)), 1,  8) -- 7597
,( 6, E,0,0,((46,49),(30,33),( 0, 1),(10,13),( 6, 9),(99,99)), 1,  8) -- 7598
,( 6, E,0,0,((48,51),(32,35),( 2, 3),(12,15),( 8,11),(99,99)), 1,  8) -- 7599
,( 6, E,0,0,((50,53),(34,37),( 4, 5),(14,17),(10,13),(99,99)), 1,  8) -- 7600
,( 6, E,0,0,((52,55),(36,39),( 6, 7),(16,19),(12,15),(99,99)), 1,  8) -- 7601
,( 6, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(16,19),(99,99)), 1,  7) -- 7602
,( 6, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(18,21),(99,99)), 1,  7) -- 7603
,( 6, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(20,23),(99,99)), 1,  7) -- 7604
,( 6, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(22,25),(99,99)), 1,  7) -- 7605
,( 6, E,0,0,((48,51),(32,35),( 0, 1),(10,13),(10,13),(99,99)), 1,  7) -- 7606
,( 6, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(12,15),(99,99)), 1,  7) -- 7607
,( 6, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(14,17),(99,99)), 1,  7) -- 7608
,( 6, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(16,19),(99,99)), 1,  7) -- 7609
,( 6, E,0,0,((50,53),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 7610
,( 6, E,0,0,((52,55),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 7611
,( 6, E,0,0,((54,57),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 7612
,( 6, E,0,0,((56,59),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 7613
,( 6, E,0,0,((50,53),(32,35),( 0, 1),(12,15),(14,17),(99,99)), 1,  7) -- 7614
,( 6, E,0,0,((52,55),(34,37),( 2, 3),(14,17),(16,19),(99,99)), 1,  7) -- 7615
,( 6, E,0,0,((54,57),(36,39),( 4, 5),(16,19),(18,21),(99,99)), 1,  7) -- 7616
,( 6, E,0,0,((56,59),(38,41),( 6, 7),(18,21),(20,23),(99,99)), 1,  7) -- 7617
,( 6, E,0,1,((50,53),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 7618
,( 6, E,0,1,((52,55),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 7619
,( 6, E,0,1,((54,57),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 7620
,( 6, E,0,1,((56,59),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 7621
,( 6, E,0,1,((50,53),(32,35),( 1, 1),(14,15),(99,99),(99,99)), 1,  7) -- 7622
,( 6, E,0,1,((52,55),(34,37),( 3, 3),(16,17),(99,99),(99,99)), 1,  7) -- 7623
,( 6, E,0,1,((54,57),(36,39),( 5, 5),(18,19),(99,99),(99,99)), 1,  7) -- 7624
,( 6, E,0,1,((56,59),(38,41),( 7, 7),(20,21),(99,99),(99,99)), 1,  7) -- 7625
,( 6, E,0,1,((46,49),(30,33),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 7626
,( 6, E,0,1,((48,51),(32,35),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 7627
,( 6, E,0,1,((50,53),(34,37),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 7628
,( 6, E,0,1,((52,55),(36,39),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 7629
,( 6, E,0,1,((50,53),(32,35),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 7630
,( 6, E,0,1,((52,55),(34,37),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 7631
,( 6, E,0,1,((54,57),(36,39),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 7632
,( 6, E,0,1,((56,59),(38,41),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 7633
,( 6, E,0,1,((54,57),(34,37),( 0, 1),(12,15),(99,99),(99,99)), 1,  6) -- 7634
,( 6, E,0,1,((56,59),(36,39),( 2, 3),(14,17),(99,99),(99,99)), 1,  6) -- 7635
,( 6, E,0,1,((58,61),(38,41),( 4, 5),(16,19),(99,99),(99,99)), 1,  6) -- 7636
,( 6, E,0,1,((60,63),(40,43),( 6, 7),(18,21),(99,99),(99,99)), 1,  6) -- 7637
,( 6, E,0,1,((42,45),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 7638
,( 6, E,0,1,((44,47),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 7639
,( 6, E,0,1,((46,49),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 7640
,( 6, E,0,1,((48,51),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 7641
,( 6, E,0,1,((54,57),(34,37),( 0, 1),( 8,11),(99,99),(99,99)), 1,  6) -- 7642
,( 6, E,0,1,((56,59),(36,39),( 2, 3),(10,13),(99,99),(99,99)), 1,  6) -- 7643
,( 6, E,0,1,((58,61),(38,41),( 4, 5),(12,15),(99,99),(99,99)), 1,  6) -- 7644
,( 6, E,0,1,((60,63),(40,43),( 6, 7),(14,17),(99,99),(99,99)), 1,  6) -- 7645
,( 6, E,0,1,((46,47),(29,29),( 0, 0),(17,17),(99,99),(99,99)), 1,  5) -- 7646
,( 6, E,0,1,((48,49),(31,31),( 2, 2),(19,19),(99,99),(99,99)), 1,  5) -- 7647
,( 6, E,0,1,((50,51),(33,33),( 4, 4),(21,21),(99,99),(99,99)), 1,  5) -- 7648
,( 6, E,0,1,((52,53),(35,35),( 6, 6),(23,23),(99,99),(99,99)), 1,  5) -- 7649
,( 6, E,0,1,((50,53),(30,31),( 0, 1),(99,99),(99,99),(99,99)), 1,  5) -- 7650
,( 6, E,0,1,((52,55),(32,33),( 2, 3),(99,99),(99,99),(99,99)), 1,  5) -- 7651
,( 6, E,0,1,((54,57),(34,35),( 4, 5),(99,99),(99,99),(99,99)), 1,  5) -- 7652
,( 6, E,0,1,((56,59),(36,37),( 6, 7),(99,99),(99,99),(99,99)), 1,  5) -- 7653
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 7654
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 7655
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 7656
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 7657
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 7658
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 7659
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 7660
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 7661
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 7662
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 7663
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 7664
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 7665
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 7666
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 7667
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 7668
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 7669
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 7670
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 7671
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 7672
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 7673
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 7674
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 7675
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 7676
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 7677
,( 6, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 7678
,( 6, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 7679
,( 6, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 7680
,( 6, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 7681
,( 6, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 7682
,( 6, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 7683
,( 6, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 7684
,( 6, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 7685
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 7686
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 7687
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 7688
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 7689
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 7690
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 7691
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 7692
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 7693
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 30) -- 7694
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 30) -- 7695
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 30) -- 7696
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 30) -- 7697
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 30) -- 7698
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 30) -- 7699
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 30) -- 7700
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 30) -- 7701
,( 6, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 30) -- 7702
,( 6, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 30) -- 7703
,( 6, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 30) -- 7704
,( 6, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 30) -- 7705
,( 6, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 30) -- 7706
,( 6, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 30) -- 7707
,( 6, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 30) -- 7708
,( 6, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 30) -- 7709
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 27) -- 7710
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 27) -- 7711
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 27) -- 7712
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 27) -- 7713
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 27) -- 7714
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 27) -- 7715
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 27) -- 7716
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 27) -- 7717
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 25) -- 7718
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 25) -- 7719
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 25) -- 7720
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 25) -- 7721
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 25) -- 7722
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 25) -- 7723
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 25) -- 7724
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 25) -- 7725
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 24) -- 7726
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 24) -- 7727
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 24) -- 7728
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 24) -- 7729
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 24) -- 7730
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 24) -- 7731
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 24) -- 7732
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 24) -- 7733
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 24) -- 7734
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 24) -- 7735
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 24) -- 7736
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 24) -- 7737
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 24) -- 7738
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 24) -- 7739
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 24) -- 7740
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 24) -- 7741
,( 6, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 23) -- 7742
,( 6, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 23) -- 7743
,( 6, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 23) -- 7744
,( 6, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 23) -- 7745
,( 6, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 23) -- 7746
,( 6, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 23) -- 7747
,( 6, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 23) -- 7748
,( 6, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 23) -- 7749
,( 6, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 23) -- 7750
,( 6, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 23) -- 7751
,( 6, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 23) -- 7752
,( 6, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 23) -- 7753
,( 6, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 23) -- 7754
,( 6, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 23) -- 7755
,( 6, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 23) -- 7756
,( 6, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 23) -- 7757
,( 6, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 22) -- 7758
,( 6, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 22) -- 7759
,( 6, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 22) -- 7760
,( 6, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 22) -- 7761
,( 6, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 22) -- 7762
,( 6, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 22) -- 7763
,( 6, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 22) -- 7764
,( 6, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 22) -- 7765
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 21) -- 7766
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 21) -- 7767
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 21) -- 7768
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 21) -- 7769
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 21) -- 7770
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 21) -- 7771
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 21) -- 7772
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 21) -- 7773
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 7774
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 7775
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 7776
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 7777
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 7778
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 7779
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 7780
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 7781
,( 6, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 20) -- 7782
,( 6, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 20) -- 7783
,( 6, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 20) -- 7784
,( 6, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 20) -- 7785
,( 6, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 20) -- 7786
,( 6, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 20) -- 7787
,( 6, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 20) -- 7788
,( 6, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 20) -- 7789
,( 6, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 20) -- 7790
,( 6, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 20) -- 7791
,( 6, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 20) -- 7792
,( 6, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 20) -- 7793
,( 6, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 20) -- 7794
,( 6, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 20) -- 7795
,( 6, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 20) -- 7796
,( 6, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 20) -- 7797
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(17,17),(10,10)), 0, 20) -- 7798
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(18,18),(11,11)), 0, 20) -- 7799
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(19,19),(12,12)), 0, 20) -- 7800
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(20,20),(13,13)), 0, 20) -- 7801
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(21,21),(14,14)), 0, 20) -- 7802
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(22,22),(15,15)), 0, 20) -- 7803
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(23,23),(16,16)), 0, 20) -- 7804
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(24,24),(17,17)), 0, 20) -- 7805
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 7806
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 7807
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 7808
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 7809
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 7810
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 7811
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 7812
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 7813
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 19) -- 7814
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 19) -- 7815
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 19) -- 7816
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 19) -- 7817
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 19) -- 7818
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 19) -- 7819
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 19) -- 7820
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 19) -- 7821
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 7822
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 7823
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 7824
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 7825
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 7826
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 7827
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 7828
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 7829
,( 6, E,0,0,((31,31),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 18) -- 7830
,( 6, E,0,0,((32,32),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 18) -- 7831
,( 6, E,0,0,((33,33),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 18) -- 7832
,( 6, E,0,0,((34,34),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 18) -- 7833
,( 6, E,0,0,((35,35),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 18) -- 7834
,( 6, E,0,0,((36,36),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 18) -- 7835
,( 6, E,0,0,((37,37),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 18) -- 7836
,( 6, E,0,0,((38,38),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 18) -- 7837
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 7838
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 7839
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 7840
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 7841
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 7842
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 7843
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 7844
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 7845
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 7846
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 7847
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 7848
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 7849
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 7850
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 7851
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 7852
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 7853
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 17) -- 7854
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 17) -- 7855
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 17) -- 7856
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 17) -- 7857
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 17) -- 7858
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 17) -- 7859
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 17) -- 7860
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 17) -- 7861
,( 6, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(11,11)), 0, 17) -- 7862
,( 6, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(12,12)), 0, 17) -- 7863
,( 6, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(13,13)), 0, 17) -- 7864
,( 6, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(14,14)), 0, 17) -- 7865
,( 6, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(15,15)), 0, 17) -- 7866
,( 6, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(16,16)), 0, 17) -- 7867
,( 6, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(17,17)), 0, 17) -- 7868
,( 6, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(18,18)), 0, 17) -- 7869
,( 6, E,0,0,((30,30),(99,99),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 7870
,( 6, E,0,0,((31,31),(99,99),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 7871
,( 6, E,0,0,((32,32),(99,99),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 7872
,( 6, E,0,0,((33,33),(99,99),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 7873
,( 6, E,0,0,((34,34),(99,99),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 7874
,( 6, E,0,0,((35,35),(99,99),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 7875
,( 6, E,0,0,((36,36),(99,99),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 7876
,( 6, E,0,0,((37,37),(99,99),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 7877
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 7878
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 7879
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 7880
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 7881
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 7882
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 7883
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 7884
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 7885
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 7886
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 7887
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 7888
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 7889
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 7890
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 7891
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 7892
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 7893
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 16) -- 7894
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 16) -- 7895
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 16) -- 7896
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 16) -- 7897
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 16) -- 7898
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 16) -- 7899
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 16) -- 7900
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 16) -- 7901
,( 6, E,0,0,((30,30),(99,99),( 0, 0),(17,17),(18,18),(12,12)), 0, 16) -- 7902
,( 6, E,0,0,((31,31),(99,99),( 1, 1),(18,18),(19,19),(13,13)), 0, 16) -- 7903
,( 6, E,0,0,((32,32),(99,99),( 2, 2),(19,19),(20,20),(14,14)), 0, 16) -- 7904
,( 6, E,0,0,((33,33),(99,99),( 3, 3),(20,20),(21,21),(15,15)), 0, 16) -- 7905
,( 6, E,0,0,((34,34),(99,99),( 4, 4),(21,21),(22,22),(16,16)), 0, 16) -- 7906
,( 6, E,0,0,((35,35),(99,99),( 5, 5),(22,22),(23,23),(17,17)), 0, 16) -- 7907
,( 6, E,0,0,((36,36),(99,99),( 6, 6),(23,23),(24,24),(18,18)), 0, 16) -- 7908
,( 6, E,0,0,((37,37),(99,99),( 7, 7),(24,24),(25,25),(19,19)), 0, 16) -- 7909
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 7910
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 7911
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 7912
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 7913
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 7914
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 7915
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 7916
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 7917
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 15) -- 7918
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 15) -- 7919
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 15) -- 7920
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 15) -- 7921
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 15) -- 7922
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 15) -- 7923
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 15) -- 7924
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 15) -- 7925
,( 6, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(12,12)), 0, 15) -- 7926
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(13,13)), 0, 15) -- 7927
,( 6, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(14,14)), 0, 15) -- 7928
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(15,15)), 0, 15) -- 7929
,( 6, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(16,16)), 0, 15) -- 7930
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(17,17)), 0, 15) -- 7931
,( 6, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(18,18)), 0, 15) -- 7932
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(19,19)), 0, 15) -- 7933
,( 6, E,0,0,((28,31),(23,23),( 0, 0),(17,17),(18,19),(10,13)), 0, 14) -- 7934
,( 6, E,0,0,((30,33),(25,25),( 2, 2),(19,19),(20,21),(12,15)), 0, 14) -- 7935
,( 6, E,0,0,((32,35),(27,27),( 4, 4),(21,21),(22,23),(14,17)), 0, 14) -- 7936
,( 6, E,0,0,((34,37),(29,29),( 6, 6),(23,23),(24,25),(16,19)), 0, 14) -- 7937
,( 6, E,0,0,((28,31),(23,23),( 0, 1),(16,17),(18,19),( 8, 9)), 0, 14) -- 7938
,( 6, E,0,0,((30,33),(25,25),( 2, 3),(18,19),(20,21),(10,11)), 0, 14) -- 7939
,( 6, E,0,0,((32,35),(27,27),( 4, 5),(20,21),(22,23),(12,13)), 0, 14) -- 7940
,( 6, E,0,0,((34,37),(29,29),( 6, 7),(22,23),(24,25),(14,15)), 0, 14) -- 7941
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(18,19),(10,11)), 0, 14) -- 7942
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(20,21),(12,13)), 0, 14) -- 7943
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(22,23),(14,15)), 0, 14) -- 7944
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(24,25),(16,17)), 0, 14) -- 7945
,( 6, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,15)), 0, 13) -- 7946
,( 6, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,17)), 0, 13) -- 7947
,( 6, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,19)), 0, 13) -- 7948
,( 6, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,21)), 0, 13) -- 7949
,( 6, E,0,0,((26,29),(99,99),( 0, 1),(18,18),(20,21),(10,13)), 0, 12) -- 7950
,( 6, E,0,0,((28,31),(99,99),( 2, 3),(20,20),(22,23),(12,15)), 0, 12) -- 7951
,( 6, E,0,0,((30,33),(99,99),( 4, 5),(22,22),(24,25),(14,17)), 0, 12) -- 7952
,( 6, E,0,0,((32,35),(99,99),( 6, 7),(24,24),(26,27),(16,19)), 0, 12) -- 7953
,( 6, E,0,0,((27,27),(99,99),( 0, 0),(17,17),(19,19),( 8,11)), 0, 12) -- 7954
,( 6, E,0,0,((29,29),(99,99),( 2, 2),(19,19),(21,21),(10,13)), 0, 12) -- 7955
,( 6, E,0,0,((31,31),(99,99),( 4, 4),(21,21),(23,23),(12,15)), 0, 12) -- 7956
,( 6, E,0,0,((33,33),(99,99),( 6, 6),(23,23),(25,25),(14,17)), 0, 12) -- 7957
,( 6, E,0,0,((27,27),(99,99),( 0, 0),(17,17),(20,20),(12,12)), 0, 12) -- 7958
,( 6, E,0,0,((29,29),(99,99),( 2, 2),(19,19),(22,22),(14,14)), 0, 12) -- 7959
,( 6, E,0,0,((31,31),(99,99),( 4, 4),(21,21),(24,24),(16,16)), 0, 12) -- 7960
,( 6, E,0,0,((33,33),(99,99),( 6, 6),(23,23),(26,26),(18,18)), 0, 12) -- 7961
,( 6, E,0,0,((28,28),(99,99),( 1, 1),(19,19),(21,21),(14,14)), 0, 12) -- 7962
,( 6, E,0,0,((30,30),(99,99),( 3, 3),(21,21),(23,23),(16,16)), 0, 12) -- 7963
,( 6, E,0,0,((32,32),(99,99),( 5, 5),(23,23),(25,25),(18,18)), 0, 12) -- 7964
,( 6, E,0,0,((34,34),(99,99),( 7, 7),(25,25),(27,27),(20,20)), 0, 12) -- 7965
,( 6, E,0,0,((27,27),(99,99),( 1, 1),(19,19),(22,22),(14,14)), 0, 12) -- 7966
,( 6, E,0,0,((29,29),(99,99),( 3, 3),(21,21),(24,24),(16,16)), 0, 12) -- 7967
,( 6, E,0,0,((31,31),(99,99),( 5, 5),(23,23),(26,26),(18,18)), 0, 12) -- 7968
,( 6, E,0,0,((33,33),(99,99),( 7, 7),(25,25),(28,28),(20,20)), 0, 12) -- 7969
,( 6, E,0,0,((26,29),(99,99),( 1, 1),(18,19),(22,22),(12,15)), 0, 11) -- 7970
,( 6, E,0,0,((28,31),(99,99),( 3, 3),(20,21),(24,24),(14,17)), 0, 11) -- 7971
,( 6, E,0,0,((30,33),(99,99),( 5, 5),(22,23),(26,26),(16,19)), 0, 11) -- 7972
,( 6, E,0,0,((32,35),(99,99),( 7, 7),(24,25),(28,28),(18,21)), 0, 11) -- 7973
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,18),(20,21),(12,15)), 0, 11) -- 7974
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,20),(22,23),(14,17)), 0, 11) -- 7975
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,22),(24,25),(16,19)), 0, 11) -- 7976
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,24),(26,27),(18,21)), 0, 11) -- 7977
,( 6, E,0,0,((24,27),(99,99),( 0, 0),(17,17),(20,21),(12,15)), 0, 11) -- 7978
,( 6, E,0,0,((26,29),(99,99),( 2, 2),(19,19),(22,23),(14,17)), 0, 11) -- 7979
,( 6, E,0,0,((28,31),(99,99),( 4, 4),(21,21),(24,25),(16,19)), 0, 11) -- 7980
,( 6, E,0,0,((30,33),(99,99),( 6, 6),(23,23),(26,27),(18,21)), 0, 11) -- 7981
,( 6, E,0,0,((28,28),(99,99),( 1, 1),(19,19),(21,21),(12,15)), 0, 11) -- 7982
,( 6, E,0,0,((30,30),(99,99),( 3, 3),(21,21),(23,23),(14,17)), 0, 11) -- 7983
,( 6, E,0,0,((32,32),(99,99),( 5, 5),(23,23),(25,25),(16,19)), 0, 11) -- 7984
,( 6, E,0,0,((34,34),(99,99),( 7, 7),(25,25),(27,27),(18,21)), 0, 11) -- 7985
,( 6, E,0,0,((26,27),(99,99),( 0, 0),(17,17),(19,19),( 7, 7)), 0, 11) -- 7986
,( 6, E,0,0,((28,29),(99,99),( 2, 2),(19,19),(21,21),( 9, 9)), 0, 11) -- 7987
,( 6, E,0,0,((30,31),(99,99),( 4, 4),(21,21),(23,23),(11,11)), 0, 11) -- 7988
,( 6, E,0,0,((32,33),(99,99),( 6, 6),(23,23),(25,25),(13,13)), 0, 11) -- 7989
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,19),(22,23),(14,17)), 0, 10) -- 7990
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,21),(24,25),(16,19)), 0, 10) -- 7991
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,23),(26,27),(18,21)), 0, 10) -- 7992
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,25),(28,29),(20,23)), 0, 10) -- 7993
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,19),(21,21),(10,13)), 0, 10) -- 7994
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,21),(23,23),(12,15)), 0, 10) -- 7995
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,23),(25,25),(14,17)), 0, 10) -- 7996
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,25),(27,27),(16,19)), 0, 10) -- 7997
,( 6, E,0,0,((26,29),(99,99),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 7998
,( 6, E,0,0,((28,31),(99,99),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 7999
,( 6, E,0,0,((30,33),(99,99),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 8000
,( 6, E,0,0,((32,35),(99,99),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 8001
,( 6, E,0,0,((26,29),(99,99),( 0, 1),(18,19),(18,19),( 6, 9)), 0, 10) -- 8002
,( 6, E,0,0,((28,31),(99,99),( 2, 3),(20,21),(20,21),( 8,11)), 0, 10) -- 8003
,( 6, E,0,0,((30,33),(99,99),( 4, 5),(22,23),(22,23),(10,13)), 0, 10) -- 8004
,( 6, E,0,0,((32,35),(99,99),( 6, 7),(24,25),(24,25),(12,15)), 0, 10) -- 8005
,( 6, E,0,0,((26,27),(99,99),( 1, 1),(20,20),(23,23),(14,17)), 0, 10) -- 8006
,( 6, E,0,0,((28,29),(99,99),( 3, 3),(22,22),(25,25),(16,19)), 0, 10) -- 8007
,( 6, E,0,0,((30,31),(99,99),( 5, 5),(24,24),(27,27),(18,21)), 0, 10) -- 8008
,( 6, E,0,0,((32,33),(99,99),( 7, 7),(26,26),(29,29),(20,23)), 0, 10) -- 8009
,( 6, E,0,0,((24,27),(99,99),( 0, 0),(17,17),(18,19),( 6, 9)), 0, 10) -- 8010
,( 6, E,0,0,((26,29),(99,99),( 2, 2),(19,19),(20,21),( 8,11)), 0, 10) -- 8011
,( 6, E,0,0,((28,31),(99,99),( 4, 4),(21,21),(22,23),(10,13)), 0, 10) -- 8012
,( 6, E,0,0,((30,33),(99,99),( 6, 6),(23,23),(24,25),(12,15)), 0, 10) -- 8013
,( 6, E,0,0,((24,27),(99,99),( 1, 1),(19,19),(22,22),(10,13)), 0, 10) -- 8014
,( 6, E,0,0,((26,29),(99,99),( 3, 3),(21,21),(24,24),(12,15)), 0, 10) -- 8015
,( 6, E,0,0,((28,31),(99,99),( 5, 5),(23,23),(26,26),(14,17)), 0, 10) -- 8016
,( 6, E,0,0,((30,33),(99,99),( 7, 7),(25,25),(28,28),(16,19)), 0, 10) -- 8017
,( 6, E,0,0,((28,28),(99,99),( 1, 1),(19,19),(20,20),(10,13)), 0, 10) -- 8018
,( 6, E,0,0,((30,30),(99,99),( 3, 3),(21,21),(22,22),(12,15)), 0, 10) -- 8019
,( 6, E,0,0,((32,32),(99,99),( 5, 5),(23,23),(24,24),(14,17)), 0, 10) -- 8020
,( 6, E,0,0,((34,34),(99,99),( 7, 7),(25,25),(26,26),(16,19)), 0, 10) -- 8021
,( 6, E,0,0,((26,26),(99,99),( 0, 0),(17,17),(20,20),( 6, 6)), 0, 10) -- 8022
,( 6, E,0,0,((28,28),(99,99),( 2, 2),(19,19),(22,22),( 8, 8)), 0, 10) -- 8023
,( 6, E,0,0,((30,30),(99,99),( 4, 4),(21,21),(24,24),(10,10)), 0, 10) -- 8024
,( 6, E,0,0,((32,32),(99,99),( 6, 6),(23,23),(26,26),(12,12)), 0, 10) -- 8025
,( 6, E,0,0,((24,24),(99,99),( 0, 0),(18,19),(23,23),(18,19)), 0, 10) -- 8026
,( 6, E,0,0,((26,26),(99,99),( 2, 2),(20,21),(25,25),(20,21)), 0, 10) -- 8027
,( 6, E,0,0,((28,28),(99,99),( 4, 4),(22,23),(27,27),(22,23)), 0, 10) -- 8028
,( 6, E,0,0,((26,26),(99,99),( 0, 0),(17,17),(20,20),(10,11)), 0, 10) -- 8029
,( 6, E,0,0,((28,28),(99,99),( 2, 2),(19,19),(22,22),(12,13)), 0, 10) -- 8030
,( 6, E,0,0,((30,30),(99,99),( 4, 4),(21,21),(24,24),(14,15)), 0, 10) -- 8031
,( 6, E,0,0,((32,32),(99,99),( 6, 6),(23,23),(26,26),(16,17)), 0, 10) -- 8032
,( 6, E,0,0,((27,27),(99,99),( 0, 0),(17,17),(17,17),( 4, 7)), 0, 10) -- 8033
,( 6, E,0,0,((29,29),(99,99),( 2, 2),(19,19),(19,19),( 6, 9)), 0, 10) -- 8034
,( 6, E,0,0,((31,31),(99,99),( 4, 4),(21,21),(21,21),( 8,11)), 0, 10) -- 8035
,( 6, E,0,0,((33,33),(99,99),( 6, 6),(23,23),(23,23),(10,13)), 0, 10) -- 8036
,( 6, E,0,0,((22,25),(99,99),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 8037
,( 6, E,0,0,((24,27),(99,99),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 8038
,( 6, E,0,0,((26,29),(99,99),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 8039
,( 6, E,0,0,((28,31),(99,99),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 8040
,( 6, E,0,0,((22,25),(99,99),( 0, 1),(18,19),(18,19),( 4, 7)), 0,  9) -- 8041
,( 6, E,0,0,((24,27),(99,99),( 2, 3),(20,21),(20,21),( 6, 9)), 0,  9) -- 8042
,( 6, E,0,0,((26,29),(99,99),( 4, 5),(22,23),(22,23),( 8,11)), 0,  9) -- 8043
,( 6, E,0,0,((28,31),(99,99),( 6, 7),(24,25),(24,25),(10,13)), 0,  9) -- 8044
,( 6, E,0,0,((24,27),(99,99),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 8045
,( 6, E,0,0,((26,29),(99,99),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 8046
,( 6, E,0,0,((28,31),(99,99),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 8047
,( 6, E,0,0,((30,33),(99,99),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 8048
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 8049
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 8050
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 8051
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 8052
,( 6, E,0,0,((22,25),(99,99),( 0, 1),(19,19),(22,23),( 8,11)), 0,  9) -- 8053
,( 6, E,0,0,((24,27),(99,99),( 2, 3),(21,21),(24,25),(10,13)), 0,  9) -- 8054
,( 6, E,0,0,((26,29),(99,99),( 4, 5),(23,23),(26,27),(12,15)), 0,  9) -- 8055
,( 6, E,0,0,((28,31),(99,99),( 6, 7),(25,25),(28,29),(14,17)), 0,  9) -- 8056
,( 6, E,0,0,((20,23),(99,99),( 0, 1),(18,19),(22,23),(12,15)), 0,  9) -- 8057
,( 6, E,0,0,((22,25),(99,99),( 2, 3),(20,21),(24,25),(14,17)), 0,  9) -- 8058
,( 6, E,0,0,((24,27),(99,99),( 4, 5),(22,23),(26,27),(16,19)), 0,  9) -- 8059
,( 6, E,0,0,((26,29),(99,99),( 6, 7),(24,25),(28,29),(18,21)), 0,  9) -- 8060
,( 6, E,0,0,((22,25),(99,99),( 0, 1),(20,21),(24,25),(14,17)), 0,  9) -- 8061
,( 6, E,0,0,((24,27),(99,99),( 2, 3),(22,23),(26,27),(16,19)), 0,  9) -- 8062
,( 6, E,0,0,((26,29),(99,99),( 4, 5),(24,25),(28,29),(18,21)), 0,  9) -- 8063
,( 6, E,0,0,((28,31),(99,99),( 6, 7),(26,27),(30,31),(20,23)), 0,  9) -- 8064
,( 6, E,0,0,((22,25),(99,99),( 1, 1),(20,20),(23,23),(15,15)), 0,  9) -- 8065
,( 6, E,0,0,((24,27),(99,99),( 3, 3),(22,22),(25,25),(17,17)), 0,  9) -- 8066
,( 6, E,0,0,((26,29),(99,99),( 5, 5),(24,24),(27,27),(19,19)), 0,  9) -- 8067
,( 6, E,0,0,((28,31),(99,99),( 7, 7),(26,26),(29,29),(21,21)), 0,  9) -- 8068
,( 6, E,0,0,((24,27),(99,99),( 0, 0),(17,17),(16,17),( 2, 2)), 0,  9) -- 8069
,( 6, E,0,0,((26,29),(99,99),( 2, 2),(19,19),(18,19),( 4, 4)), 0,  9) -- 8070
,( 6, E,0,0,((28,31),(99,99),( 4, 4),(21,21),(20,21),( 6, 6)), 0,  9) -- 8071
,( 6, E,0,0,((30,33),(99,99),( 6, 6),(23,23),(22,23),( 8, 8)), 0,  9) -- 8072
,( 6, E,0,0,((22,25),(99,99),( 0, 1),(18,18),(20,21),(10,11)), 0,  9) -- 8073
,( 6, E,0,0,((24,27),(99,99),( 2, 3),(20,20),(22,23),(12,13)), 0,  9) -- 8074
,( 6, E,0,0,((26,29),(99,99),( 4, 5),(22,22),(24,25),(14,15)), 0,  9) -- 8075
,( 6, E,0,0,((28,31),(99,99),( 6, 7),(24,24),(26,27),(16,17)), 0,  9) -- 8076
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(19,19),(22,22),( 6, 9)), 0,  9) -- 8077
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(21,21),(24,24),( 8,11)), 0,  9) -- 8078
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(23,23),(26,26),(10,13)), 0,  9) -- 8079
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(25,25),(28,28),(12,15)), 0,  9) -- 8080
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,19),(20,21),( 0, 1)), 0,  9) -- 8081
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,21),(22,23),( 2, 3)), 0,  9) -- 8082
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,23),(24,25),( 4, 5)), 0,  9) -- 8083
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,25),(26,27),( 6, 7)), 0,  9) -- 8084
,( 6, E,0,0,((24,27),(99,99),( 0, 0),(17,17),(18,19),( 2, 5)), 0,  9) -- 8085
,( 6, E,0,0,((26,29),(99,99),( 2, 2),(19,19),(20,21),( 4, 7)), 0,  9) -- 8086
,( 6, E,0,0,((28,31),(99,99),( 4, 4),(21,21),(22,23),( 6, 9)), 0,  9) -- 8087
,( 6, E,0,0,((30,33),(99,99),( 6, 6),(23,23),(24,25),( 8,11)), 0,  9) -- 8088
,( 6, E,0,0,((22,25),(99,99),( 0, 0),(18,18),(18,19),( 0, 3)), 0,  9) -- 8089
,( 6, E,0,0,((24,27),(99,99),( 2, 2),(20,20),(20,21),( 2, 5)), 0,  9) -- 8090
,( 6, E,0,0,((26,29),(99,99),( 4, 4),(22,22),(22,23),( 4, 7)), 0,  9) -- 8091
,( 6, E,0,0,((28,31),(99,99),( 6, 6),(24,24),(24,25),( 6, 9)), 0,  9) -- 8092
,( 6, E,0,0,((24,27),(99,99),( 1, 1),(20,20),(22,23),( 6, 9)), 0,  9) -- 8093
,( 6, E,0,0,((26,29),(99,99),( 3, 3),(22,22),(24,25),( 8,11)), 0,  9) -- 8094
,( 6, E,0,0,((28,31),(99,99),( 5, 5),(24,24),(26,27),(10,13)), 0,  9) -- 8095
,( 6, E,0,0,((30,33),(99,99),( 7, 7),(26,26),(28,29),(12,15)), 0,  9) -- 8096
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,19),(16,17),(99,99)), 0,  9) -- 8097
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,21),(18,19),(99,99)), 0,  9) -- 8098
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,23),(20,21),(99,99)), 0,  9) -- 8099
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,25),(22,23),(99,99)), 0,  9) -- 8100
,( 6, E,0,0,((20,23),(99,99),( 0, 1),(18,21),(20,23),(12,12)), 0,  8) -- 8101
,( 6, E,0,0,((22,25),(99,99),( 2, 3),(20,23),(22,25),(14,14)), 0,  8) -- 8102
,( 6, E,0,0,((24,27),(99,99),( 4, 5),(22,25),(24,27),(16,16)), 0,  8) -- 8103
,( 6, E,0,0,((26,29),(99,99),( 6, 7),(24,27),(26,29),(18,18)), 0,  8) -- 8104
,( 6, E,0,0,((24,27),(99,99),( 0, 1),(18,21),(20,23),(12,12)), 0,  8) -- 8105
,( 6, E,0,0,((26,29),(99,99),( 2, 3),(20,23),(22,25),(14,14)), 0,  8) -- 8106
,( 6, E,0,0,((28,31),(99,99),( 4, 5),(22,25),(24,27),(16,16)), 0,  8) -- 8107
,( 6, E,0,0,((30,33),(99,99),( 6, 7),(24,27),(26,29),(18,18)), 0,  8) -- 8108
,( 6, E,0,0,((20,23),(99,99),( 0, 1),(18,21),(16,19),(99,99)), 0,  8) -- 8109
,( 6, E,0,0,((22,25),(99,99),( 2, 3),(20,23),(18,21),(99,99)), 0,  8) -- 8110
,( 6, E,0,0,((24,27),(99,99),( 4, 5),(22,25),(20,23),(99,99)), 0,  8) -- 8111
,( 6, E,0,0,((26,29),(99,99),( 6, 7),(24,27),(22,25),(99,99)), 0,  8) -- 8112
,( 6, E,0,1,((20,23),(99,99),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 8113
,( 6, E,0,1,((22,25),(99,99),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 8114
,( 6, E,0,1,((24,27),(99,99),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 8115
,( 6, E,0,1,((26,29),(99,99),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 8116
,( 6, E,0,1,((16,19),(99,99),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 8117
,( 6, E,0,1,((18,21),(99,99),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 8118
,( 6, E,0,1,((20,23),(99,99),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 8119
,( 6, E,0,1,((22,25),(99,99),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 8120
,( 6, E,0,1,((22,25),(99,99),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 8121
,( 6, E,0,1,((24,27),(99,99),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 8122
,( 6, E,0,1,((26,29),(99,99),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 8123
,( 6, E,0,1,((28,31),(99,99),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 8124
,( 6, E,0,1,((18,21),(99,99),( 0, 1),(16,17),(99,99),(99,99)), 0,  7) -- 8125
,( 6, E,0,1,((20,23),(99,99),( 2, 3),(18,19),(99,99),(99,99)), 0,  7) -- 8126
,( 6, E,0,1,((22,25),(99,99),( 4, 5),(20,21),(99,99),(99,99)), 0,  7) -- 8127
,( 6, E,0,1,((24,27),(99,99),( 6, 7),(22,23),(99,99),(99,99)), 0,  7) -- 8128
,( 6, E,0,1,((14,17),(99,99),( 0, 1),(20,23),(99,99),(99,99)), 0,  7) -- 8129
,( 6, E,0,1,((16,19),(99,99),( 2, 3),(22,25),(99,99),(99,99)), 0,  7) -- 8130
,( 6, E,0,1,((18,21),(99,99),( 4, 5),(24,27),(99,99),(99,99)), 0,  7) -- 8131
,( 6, E,0,1,((20,23),(99,99),( 6, 7),(26,29),(99,99),(99,99)), 0,  7) -- 8132
,( 6, E,0,1,((22,25),(99,99),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 8133
,( 6, E,0,1,((24,27),(99,99),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 8134
,( 6, E,0,1,((26,29),(99,99),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 8135
,( 6, E,0,1,((28,31),(99,99),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 8136
,( 6, E,0,1,((12,15),(99,99),( 0, 1),(18,21),(99,99),(99,99)), 0,  6) -- 8137
,( 6, E,0,1,((14,17),(99,99),( 2, 3),(20,23),(99,99),(99,99)), 0,  6) -- 8138
,( 6, E,0,1,((16,19),(99,99),( 4, 5),(22,25),(99,99),(99,99)), 0,  6) -- 8139
,( 6, E,0,1,((18,21),(99,99),( 6, 7),(24,27),(99,99),(99,99)), 0,  6) -- 8140
,( 6, E,0,1,((26,29),(99,99),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 8141
,( 6, E,0,1,((28,31),(99,99),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 8142
,( 6, E,0,1,((30,33),(99,99),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 8143
,( 6, E,0,1,((32,35),(99,99),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 8144
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 31) -- 8145
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 31) -- 8146
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 1, 31) -- 8147
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 1, 31) -- 8148
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 1, 31) -- 8149
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 1, 31) -- 8150
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 1, 31) -- 8151
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 1, 31) -- 8152
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 8153
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 8154
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 8155
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 8156
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 8157
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 8158
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 8159
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 8160
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 8161
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 8162
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 8163
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 8164
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 8165
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 8166
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 8167
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 8168
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 8169
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 8170
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 8171
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 8172
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 8173
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 8174
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 8175
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 8176
,( 7, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 8177
,( 7, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 8178
,( 7, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 8179
,( 7, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 8180
,( 7, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 8181
,( 7, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 8182
,( 7, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 8183
,( 7, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 8184
,( 7, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 8185
,( 7, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 8186
,( 7, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 8187
,( 7, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 8188
,( 7, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 8189
,( 7, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 8190
,( 7, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 8191
,( 7, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 8192
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 1, 31) -- 8193
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 1, 31) -- 8194
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 1, 31) -- 8195
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 1, 31) -- 8196
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 1, 31) -- 8197
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 1, 31) -- 8198
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 1, 31) -- 8199
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 1, 31) -- 8200
,( 7, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 8201
,( 7, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 8202
,( 7, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 8203
,( 7, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 8204
,( 7, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 8205
,( 7, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 8206
,( 7, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 8207
,( 7, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 8208
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 30) -- 8209
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 30) -- 8210
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 30) -- 8211
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 30) -- 8212
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 30) -- 8213
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 30) -- 8214
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 30) -- 8215
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 30) -- 8216
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 28) -- 8217
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 28) -- 8218
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 28) -- 8219
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 28) -- 8220
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 28) -- 8221
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 28) -- 8222
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 28) -- 8223
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 28) -- 8224
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 27) -- 8225
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 27) -- 8226
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 27) -- 8227
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 27) -- 8228
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 27) -- 8229
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 27) -- 8230
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 27) -- 8231
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 27) -- 8232
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 26) -- 8233
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 26) -- 8234
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 26) -- 8235
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 26) -- 8236
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 26) -- 8237
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 26) -- 8238
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 26) -- 8239
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 26) -- 8240
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 25) -- 8241
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 25) -- 8242
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 25) -- 8243
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 25) -- 8244
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 25) -- 8245
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 25) -- 8246
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 25) -- 8247
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 25) -- 8248
,( 7, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 8249
,( 7, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 8250
,( 7, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 8251
,( 7, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 8252
,( 7, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 8253
,( 7, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 8254
,( 7, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 8255
,( 7, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 8256
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 23) -- 8257
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 23) -- 8258
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 23) -- 8259
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 23) -- 8260
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 23) -- 8261
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 23) -- 8262
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 23) -- 8263
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 23) -- 8264
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 23) -- 8265
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 23) -- 8266
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 23) -- 8267
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 23) -- 8268
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 23) -- 8269
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 23) -- 8270
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 23) -- 8271
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 23) -- 8272
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 8273
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 8274
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 8275
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 8276
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 8277
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 8278
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 8279
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 8280
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 22) -- 8281
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 22) -- 8282
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),(10,10)), 1, 22) -- 8283
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(11,11)), 1, 22) -- 8284
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(12,12)), 1, 22) -- 8285
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(13,13)), 1, 22) -- 8286
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(14,14)), 1, 22) -- 8287
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(15,15)), 1, 22) -- 8288
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 21) -- 8289
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 21) -- 8290
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 21) -- 8291
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 21) -- 8292
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 21) -- 8293
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 21) -- 8294
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 21) -- 8295
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 21) -- 8296
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 21) -- 8297
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 21) -- 8298
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 21) -- 8299
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 21) -- 8300
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 21) -- 8301
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 21) -- 8302
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 21) -- 8303
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 21) -- 8304
,( 7, E,0,0,((33,33),(26,26),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 20) -- 8305
,( 7, E,0,0,((34,34),(27,27),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 20) -- 8306
,( 7, E,0,0,((35,35),(28,28),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 20) -- 8307
,( 7, E,0,0,((36,36),(29,29),( 3, 3),(19,19),(19,19),(10,10)), 1, 20) -- 8308
,( 7, E,0,0,((37,37),(30,30),( 4, 4),(20,20),(20,20),(11,11)), 1, 20) -- 8309
,( 7, E,0,0,((38,38),(31,31),( 5, 5),(21,21),(21,21),(12,12)), 1, 20) -- 8310
,( 7, E,0,0,((39,39),(32,32),( 6, 6),(22,22),(22,22),(13,13)), 1, 20) -- 8311
,( 7, E,0,0,((40,40),(33,33),( 7, 7),(23,23),(23,23),(14,14)), 1, 20) -- 8312
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 19) -- 8313
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 19) -- 8314
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 19) -- 8315
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(19,19),(19,19),(10,10)), 1, 19) -- 8316
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(20,20),(20,20),(11,11)), 1, 19) -- 8317
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(21,21),(21,21),(12,12)), 1, 19) -- 8318
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(22,22),(22,22),(13,13)), 1, 19) -- 8319
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(23,23),(23,23),(14,14)), 1, 19) -- 8320
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 19) -- 8321
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 19) -- 8322
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 19) -- 8323
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(19,19),(10,10)), 1, 19) -- 8324
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(20,20),(11,11)), 1, 19) -- 8325
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(21,21),(12,12)), 1, 19) -- 8326
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(22,22),(13,13)), 1, 19) -- 8327
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(23,23),(14,14)), 1, 19) -- 8328
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 6, 6)), 1, 19) -- 8329
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 7, 7)), 1, 19) -- 8330
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 8, 8)), 1, 19) -- 8331
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),( 9, 9)), 1, 19) -- 8332
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(10,10)), 1, 19) -- 8333
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(11,11)), 1, 19) -- 8334
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(12,12)), 1, 19) -- 8335
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(13,13)), 1, 19) -- 8336
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 8337
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 8338
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 8339
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 8340
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 8341
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 8342
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 8343
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 8344
,( 7, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 19) -- 8345
,( 7, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 19) -- 8346
,( 7, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 19) -- 8347
,( 7, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 19) -- 8348
,( 7, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 19) -- 8349
,( 7, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(10,10)), 1, 19) -- 8350
,( 7, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(11,11)), 1, 19) -- 8351
,( 7, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(12,12)), 1, 19) -- 8352
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 8353
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 8354
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 8355
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 8356
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 8357
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 8358
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 8359
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 8360
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 8361
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 8362
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 8363
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 8364
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 8365
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 8366
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 8367
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 8368
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 18) -- 8369
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 18) -- 8370
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 18) -- 8371
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 18) -- 8372
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 18) -- 8373
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 18) -- 8374
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 18) -- 8375
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 18) -- 8376
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(16,16),( 6, 6)), 1, 18) -- 8377
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(17,17),( 7, 7)), 1, 18) -- 8378
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(18,18),( 8, 8)), 1, 18) -- 8379
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(19,19),( 9, 9)), 1, 18) -- 8380
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(20,20),(10,10)), 1, 18) -- 8381
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(21,21),(11,11)), 1, 18) -- 8382
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(22,22),(12,12)), 1, 18) -- 8383
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(23,23),(13,13)), 1, 18) -- 8384
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 8385
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 8386
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 8387
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 8388
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 8389
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 8390
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 8391
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 8392
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 8393
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 8394
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 8395
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 8396
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 8397
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 8398
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 8399
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 8400
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 8401
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 8402
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 8403
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 8404
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 8405
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 8406
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 8407
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 8408
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 8409
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 8410
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 8411
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 8412
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 8413
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 8414
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 8415
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 8416
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 17) -- 8417
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 17) -- 8418
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 17) -- 8419
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 17) -- 8420
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 17) -- 8421
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(10,10)), 1, 17) -- 8422
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(11,11)), 1, 17) -- 8423
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(12,12)), 1, 17) -- 8424
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 8425
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 8426
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 8427
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 8428
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 8429
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 8430
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 8431
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 8432
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 8433
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 8434
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 8435
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 8436
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 8437
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 8438
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 8439
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 8440
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 8441
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 8442
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 8443
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 8444
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 8445
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 8446
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 8447
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 8448
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 17) -- 8449
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 17) -- 8450
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 17) -- 8451
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 17) -- 8452
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 17) -- 8453
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 17) -- 8454
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 17) -- 8455
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 17) -- 8456
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 8457
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 8458
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 8459
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 8460
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 8461
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 8462
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 8463
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 8464
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 8465
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 8466
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 8467
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 8468
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 8469
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 8470
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 8471
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 8472
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 16) -- 8473
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 16) -- 8474
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 16) -- 8475
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 16) -- 8476
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 16) -- 8477
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(19,19),(19,19),(10,10)), 1, 16) -- 8478
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(20,20),(20,20),(11,11)), 1, 16) -- 8479
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(21,21),(21,21),(12,12)), 1, 16) -- 8480
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 8481
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 8482
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 8483
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 8484
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 8485
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 8486
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 8487
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 8488
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 16) -- 8489
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 16) -- 8490
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 16) -- 8491
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 16) -- 8492
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 16) -- 8493
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 16) -- 8494
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(20,20),(20,20),(10,10)), 1, 16) -- 8495
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(21,21),(21,21),(11,11)), 1, 16) -- 8496
,( 7, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 16) -- 8497
,( 7, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 16) -- 8498
,( 7, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 16) -- 8499
,( 7, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 16) -- 8500
,( 7, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 16) -- 8501
,( 7, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 16) -- 8502
,( 7, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(10,10)), 1, 16) -- 8503
,( 7, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(11,11)), 1, 16) -- 8504
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 15) -- 8505
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 15) -- 8506
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 15) -- 8507
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 15) -- 8508
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 15) -- 8509
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),(10,10)), 1, 15) -- 8510
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(11,11)), 1, 15) -- 8511
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(12,12)), 1, 15) -- 8512
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 8513
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 8514
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 8515
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 8516
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 8517
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 8518
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 8519
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 8520
,( 7, E,0,0,((34,34),(26,26),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 8521
,( 7, E,0,0,((35,35),(27,27),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 8522
,( 7, E,0,0,((36,36),(28,28),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 8523
,( 7, E,0,0,((37,37),(29,29),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 8524
,( 7, E,0,0,((38,38),(30,30),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 8525
,( 7, E,0,0,((39,39),(31,31),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 8526
,( 7, E,0,0,((40,40),(32,32),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 8527
,( 7, E,0,0,((41,41),(33,33),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 8528
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 15) -- 8529
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 15) -- 8530
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 15) -- 8531
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 15) -- 8532
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 15) -- 8533
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 15) -- 8534
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(10,10)), 1, 15) -- 8535
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(11,11)), 1, 15) -- 8536
,( 7, E,0,0,((36,36),(27,27),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 8537
,( 7, E,0,0,((37,37),(28,28),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 8538
,( 7, E,0,0,((38,38),(29,29),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 8539
,( 7, E,0,0,((39,39),(30,30),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 8540
,( 7, E,0,0,((40,40),(31,31),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 8541
,( 7, E,0,0,((41,41),(32,32),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 8542
,( 7, E,0,0,((42,42),(33,33),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 8543
,( 7, E,0,0,((43,43),(34,34),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 8544
,( 7, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 8545
,( 7, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 8546
,( 7, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 8547
,( 7, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 8548
,( 7, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 8549
,( 7, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 8550
,( 7, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 8551
,( 7, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 8552
,( 7, E,0,0,((35,35),(27,27),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 8553
,( 7, E,0,0,((36,36),(28,28),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 8554
,( 7, E,0,0,((37,37),(29,29),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 8555
,( 7, E,0,0,((38,38),(30,30),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 8556
,( 7, E,0,0,((39,39),(31,31),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 8557
,( 7, E,0,0,((40,40),(32,32),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 8558
,( 7, E,0,0,((41,41),(33,33),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 8559
,( 7, E,0,0,((42,42),(34,34),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 8560
,( 7, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 8561
,( 7, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 8562
,( 7, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 8563
,( 7, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 8564
,( 7, E,0,0,((36,39),(28,29),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 8565
,( 7, E,0,0,((38,41),(30,31),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 8566
,( 7, E,0,0,((40,43),(32,33),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 8567
,( 7, E,0,0,((42,45),(34,35),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 8568
,( 7, E,0,0,((34,37),(26,27),( 0, 0),(14,15),(13,13),( 2, 5)), 1, 14) -- 8569
,( 7, E,0,0,((36,39),(28,29),( 2, 2),(16,17),(15,15),( 4, 7)), 1, 14) -- 8570
,( 7, E,0,0,((38,41),(30,31),( 4, 4),(18,19),(17,17),( 6, 9)), 1, 14) -- 8571
,( 7, E,0,0,((40,43),(32,33),( 6, 6),(20,21),(19,19),( 8,11)), 1, 14) -- 8572
,( 7, E,0,0,((36,39),(28,29),( 0, 1),(15,15),(14,15),( 4, 7)), 1, 13) -- 8573
,( 7, E,0,0,((38,41),(30,31),( 2, 3),(17,17),(16,17),( 6, 9)), 1, 13) -- 8574
,( 7, E,0,0,((40,43),(32,33),( 4, 5),(19,19),(18,19),( 8,11)), 1, 13) -- 8575
,( 7, E,0,0,((42,45),(34,35),( 6, 7),(21,21),(20,21),(10,13)), 1, 13) -- 8576
,( 7, E,0,0,((36,39),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 8577
,( 7, E,0,0,((38,41),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 8578
,( 7, E,0,0,((40,43),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 8579
,( 7, E,0,0,((42,45),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 8580
,( 7, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 8581
,( 7, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 8582
,( 7, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 8583
,( 7, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 8584
,( 7, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,13),( 2, 5)), 1, 12) -- 8585
,( 7, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,15),( 4, 7)), 1, 12) -- 8586
,( 7, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,17),( 6, 9)), 1, 12) -- 8587
,( 7, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,19),( 8,11)), 1, 12) -- 8588
,( 7, E,0,0,((40,41),(29,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 8589
,( 7, E,0,0,((42,43),(31,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 8590
,( 7, E,0,0,((44,45),(33,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 8591
,( 7, E,0,0,((46,47),(35,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 8592
,( 7, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 8593
,( 7, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 8594
,( 7, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(10,13)), 1, 11) -- 8595
,( 7, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(12,15)), 1, 11) -- 8596
,( 7, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),( 2, 5)), 1, 11) -- 8597
,( 7, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),( 4, 7)), 1, 11) -- 8598
,( 7, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),( 6, 9)), 1, 11) -- 8599
,( 7, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),( 8,11)), 1, 11) -- 8600
,( 7, E,0,0,((38,41),(28,29),( 0, 1),(12,13),(10,11),( 0, 3)), 1, 11) -- 8601
,( 7, E,0,0,((40,43),(30,31),( 2, 3),(14,15),(12,13),( 2, 5)), 1, 11) -- 8602
,( 7, E,0,0,((42,45),(32,33),( 4, 5),(16,17),(14,15),( 4, 7)), 1, 11) -- 8603
,( 7, E,0,0,((44,47),(34,35),( 6, 7),(18,19),(16,17),( 6, 9)), 1, 11) -- 8604
,( 7, E,0,0,((40,43),(30,31),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 11) -- 8605
,( 7, E,0,0,((42,45),(32,33),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 11) -- 8606
,( 7, E,0,0,((44,47),(34,35),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 11) -- 8607
,( 7, E,0,0,((46,49),(36,37),( 7, 7),(20,21),(18,19),( 8,11)), 1, 11) -- 8608
,( 7, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 8609
,( 7, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 8610
,( 7, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 8611
,( 7, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 8612
,( 7, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,14),( 4, 5)), 1, 11) -- 8613
,( 7, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,16),( 6, 7)), 1, 11) -- 8614
,( 7, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,18),( 8, 9)), 1, 11) -- 8615
,( 7, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,20),(10,11)), 1, 11) -- 8616
,( 7, E,0,0,((40,43),(30,31),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 10) -- 8617
,( 7, E,0,0,((42,45),(32,33),( 2, 3),(16,17),(16,17),( 8,11)), 1, 10) -- 8618
,( 7, E,0,0,((44,47),(34,35),( 4, 5),(18,19),(18,19),(10,13)), 1, 10) -- 8619
,( 7, E,0,0,((46,49),(36,37),( 6, 7),(20,21),(20,21),(12,15)), 1, 10) -- 8620
,( 7, E,0,0,((40,43),(30,31),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 8621
,( 7, E,0,0,((42,45),(32,33),( 2, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 8622
,( 7, E,0,0,((44,47),(34,35),( 4, 5),(18,19),(16,17),(10,13)), 1, 10) -- 8623
,( 7, E,0,0,((46,49),(36,37),( 6, 7),(20,21),(18,19),(12,15)), 1, 10) -- 8624
,( 7, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(12,13),( 6, 9)), 1, 10) -- 8625
,( 7, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(14,15),( 8,11)), 1, 10) -- 8626
,( 7, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(16,17),(10,13)), 1, 10) -- 8627
,( 7, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(18,19),(12,15)), 1, 10) -- 8628
,( 7, E,0,0,((40,43),(30,31),( 0, 1),(12,13),(10,11),( 0, 3)), 1, 10) -- 8629
,( 7, E,0,0,((42,45),(32,33),( 2, 3),(14,15),(12,13),( 2, 5)), 1, 10) -- 8630
,( 7, E,0,0,((44,47),(34,35),( 4, 5),(16,17),(14,15),( 4, 7)), 1, 10) -- 8631
,( 7, E,0,0,((46,49),(36,37),( 6, 7),(18,19),(16,17),( 6, 9)), 1, 10) -- 8632
,( 7, E,0,0,((40,43),(30,31),( 1, 1),(14,14),(10,11),( 0, 3)), 1, 10) -- 8633
,( 7, E,0,0,((42,45),(32,33),( 3, 3),(16,16),(12,13),( 2, 5)), 1, 10) -- 8634
,( 7, E,0,0,((44,47),(34,35),( 5, 5),(18,18),(14,15),( 4, 7)), 1, 10) -- 8635
,( 7, E,0,0,((46,49),(36,37),( 7, 7),(20,20),(16,17),( 6, 9)), 1, 10) -- 8636
,( 7, E,0,0,((38,41),(28,29),( 0, 0),(13,13),(11,11),( 4, 7)), 1, 10) -- 8637
,( 7, E,0,0,((40,43),(30,31),( 2, 2),(15,15),(13,13),( 6, 9)), 1, 10) -- 8638
,( 7, E,0,0,((42,45),(32,33),( 4, 4),(17,17),(15,15),( 8,11)), 1, 10) -- 8639
,( 7, E,0,0,((44,47),(34,35),( 6, 6),(19,19),(17,17),(10,13)), 1, 10) -- 8640
,( 7, E,0,0,((40,41),(29,29),( 0, 1),(14,14),(11,11),( 0, 3)), 1, 10) -- 8641
,( 7, E,0,0,((42,43),(31,31),( 2, 3),(16,16),(13,13),( 2, 5)), 1, 10) -- 8642
,( 7, E,0,0,((44,45),(33,33),( 4, 5),(18,18),(15,15),( 4, 7)), 1, 10) -- 8643
,( 7, E,0,0,((46,47),(35,35),( 6, 7),(20,20),(17,17),( 6, 9)), 1, 10) -- 8644
,( 7, E,0,0,((36,39),(27,27),( 0, 0),(14,15),(14,14),( 6, 9)), 1, 10) -- 8645
,( 7, E,0,0,((38,41),(29,29),( 2, 2),(16,17),(16,16),( 8,11)), 1, 10) -- 8646
,( 7, E,0,0,((40,43),(31,31),( 4, 4),(18,19),(18,18),(10,13)), 1, 10) -- 8647
,( 7, E,0,0,((42,45),(33,33),( 6, 6),(20,21),(20,20),(12,15)), 1, 10) -- 8648
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 8649
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 8650
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 8651
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 8652
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 6, 9)), 1,  9) -- 8653
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),( 8,11)), 1,  9) -- 8654
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(10,13)), 1,  9) -- 8655
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(12,15)), 1,  9) -- 8656
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 8657
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 8658
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 8659
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 8660
,( 7, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(12,13),( 8,11)), 1,  9) -- 8661
,( 7, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(14,15),(10,13)), 1,  9) -- 8662
,( 7, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(16,17),(12,15)), 1,  9) -- 8663
,( 7, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(18,19),(14,17)), 1,  9) -- 8664
,( 7, E,0,0,((44,47),(32,33),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 8665
,( 7, E,0,0,((46,49),(34,35),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 8666
,( 7, E,0,0,((48,51),(36,37),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 8667
,( 7, E,0,0,((50,53),(38,39),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 8668
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 8669
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 8670
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 8671
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 8672
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),(10,11)), 1,  9) -- 8673
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(12,13)), 1,  9) -- 8674
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(14,15)), 1,  9) -- 8675
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(16,17)), 1,  9) -- 8676
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(12,13),( 4, 7)), 1,  9) -- 8677
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(14,15),( 6, 9)), 1,  9) -- 8678
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(16,17),( 8,11)), 1,  9) -- 8679
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(18,19),(10,13)), 1,  9) -- 8680
,( 7, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 8681
,( 7, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 8682
,( 7, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 8683
,( 7, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 8684
,( 7, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(12,13),( 8,11)), 1,  9) -- 8685
,( 7, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(14,15),(10,13)), 1,  9) -- 8686
,( 7, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(16,17),(12,15)), 1,  9) -- 8687
,( 7, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(18,19),(14,17)), 1,  9) -- 8688
,( 7, E,0,0,((44,47),(32,32),( 1, 1),(14,15),(12,13),( 6, 9)), 1,  9) -- 8689
,( 7, E,0,0,((46,49),(34,34),( 3, 3),(16,17),(14,15),( 8,11)), 1,  9) -- 8690
,( 7, E,0,0,((48,51),(36,36),( 5, 5),(18,19),(16,17),(10,13)), 1,  9) -- 8691
,( 7, E,0,0,((50,53),(38,38),( 7, 7),(20,21),(18,19),(12,15)), 1,  9) -- 8692
,( 7, E,0,0,((40,43),(30,31),( 0, 0),(12,13),(11,11),( 8, 9)), 1,  9) -- 8693
,( 7, E,0,0,((42,45),(32,33),( 2, 2),(14,15),(13,13),(10,11)), 1,  9) -- 8694
,( 7, E,0,0,((44,47),(34,35),( 4, 4),(16,17),(15,15),(12,13)), 1,  9) -- 8695
,( 7, E,0,0,((46,49),(36,37),( 6, 6),(18,19),(17,17),(14,15)), 1,  9) -- 8696
,( 7, E,0,0,((40,43),(30,31),( 0, 1),(13,13),(12,12),( 2, 5)), 1,  9) -- 8697
,( 7, E,0,0,((42,45),(32,33),( 2, 3),(15,15),(14,14),( 4, 7)), 1,  9) -- 8698
,( 7, E,0,0,((44,47),(34,35),( 4, 5),(17,17),(16,16),( 6, 9)), 1,  9) -- 8699
,( 7, E,0,0,((46,49),(36,37),( 6, 7),(19,19),(18,18),( 8,11)), 1,  9) -- 8700
,( 7, E,0,0,((44,47),(32,33),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 8701
,( 7, E,0,0,((46,49),(34,35),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 8702
,( 7, E,0,0,((48,51),(36,37),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 8703
,( 7, E,0,0,((50,53),(38,39),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 8704
,( 7, E,0,0,((40,43),(29,29),( 0, 0),(12,13),(11,11),( 4, 7)), 1,  9) -- 8705
,( 7, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(13,13),( 6, 9)), 1,  9) -- 8706
,( 7, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(15,15),( 8,11)), 1,  9) -- 8707
,( 7, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(17,17),(10,13)), 1,  9) -- 8708
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(14,15),(12,12)), 1,  9) -- 8709
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(16,17),(14,14)), 1,  9) -- 8710
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(18,19),(16,16)), 1,  9) -- 8711
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(20,21),(18,18)), 1,  9) -- 8712
,( 7, E,0,0,((40,43),(30,31),( 1, 1),(15,15),(16,16),(12,15)), 1,  9) -- 8713
,( 7, E,0,0,((42,45),(32,33),( 3, 3),(17,17),(18,18),(14,17)), 1,  9) -- 8714
,( 7, E,0,0,((44,47),(34,35),( 5, 5),(19,19),(20,20),(16,19)), 1,  9) -- 8715
,( 7, E,0,0,((46,49),(36,37),( 7, 7),(21,21),(22,22),(18,21)), 1,  9) -- 8716
,( 7, E,0,0,((41,41),(29,29),( 0, 0),(12,12),( 9, 9),( 0, 3)), 1,  9) -- 8717
,( 7, E,0,0,((43,43),(31,31),( 2, 2),(14,14),(11,11),( 2, 5)), 1,  9) -- 8718
,( 7, E,0,0,((45,45),(33,33),( 4, 4),(16,16),(13,13),( 4, 7)), 1,  9) -- 8719
,( 7, E,0,0,((47,47),(35,35),( 6, 6),(18,18),(15,15),( 6, 9)), 1,  9) -- 8720
,( 7, E,0,0,((38,41),(28,29),( 0, 0),(14,14),(13,13),(10,11)), 1,  9) -- 8721
,( 7, E,0,0,((40,43),(30,31),( 2, 2),(16,16),(15,15),(12,13)), 1,  9) -- 8722
,( 7, E,0,0,((42,45),(32,33),( 4, 4),(18,18),(17,17),(14,15)), 1,  9) -- 8723
,( 7, E,0,0,((44,47),(34,35),( 6, 6),(20,20),(19,19),(16,17)), 1,  9) -- 8724
,( 7, E,0,0,((44,47),(32,33),( 0, 1),(12,13),(12,13),( 6, 9)), 1,  9) -- 8725
,( 7, E,0,0,((46,49),(34,35),( 2, 3),(14,15),(14,15),( 8,11)), 1,  9) -- 8726
,( 7, E,0,0,((48,51),(36,37),( 4, 5),(16,17),(16,17),(10,13)), 1,  9) -- 8727
,( 7, E,0,0,((50,53),(38,39),( 6, 7),(18,19),(18,19),(12,15)), 1,  9) -- 8728
,( 7, E,0,0,((42,42),(29,29),( 0, 0),(12,13),(12,12),( 4, 7)), 1,  9) -- 8729
,( 7, E,0,0,((44,44),(31,31),( 2, 2),(14,15),(14,14),( 6, 9)), 1,  9) -- 8730
,( 7, E,0,0,((46,46),(33,33),( 4, 4),(16,17),(16,16),( 8,11)), 1,  9) -- 8731
,( 7, E,0,0,((48,48),(35,35),( 6, 6),(18,19),(18,18),(10,13)), 1,  9) -- 8732
,( 7, E,0,0,((44,45),(32,32),( 1, 1),(14,14),(10,11),( 0, 3)), 1,  9) -- 8733
,( 7, E,0,0,((46,47),(34,34),( 3, 3),(16,16),(12,13),( 2, 5)), 1,  9) -- 8734
,( 7, E,0,0,((48,49),(36,36),( 5, 5),(18,18),(14,15),( 4, 7)), 1,  9) -- 8735
,( 7, E,0,0,((50,51),(38,38),( 7, 7),(20,20),(16,17),( 6, 9)), 1,  9) -- 8736
,( 7, E,0,0,((44,47),(32,33),( 0, 1),(12,13),(10,11),( 2, 3)), 1,  9) -- 8737
,( 7, E,0,0,((46,49),(34,35),( 2, 3),(14,15),(12,13),( 4, 5)), 1,  9) -- 8738
,( 7, E,0,0,((48,51),(36,37),( 4, 5),(16,17),(14,15),( 6, 7)), 1,  9) -- 8739
,( 7, E,0,0,((50,53),(38,39),( 6, 7),(18,19),(16,17),( 8, 9)), 1,  9) -- 8740
,( 7, E,0,0,((41,41),(30,30),( 1, 1),(14,15),(14,14),(10,13)), 1,  9) -- 8741
,( 7, E,0,0,((43,43),(32,32),( 3, 3),(16,17),(16,16),(12,15)), 1,  9) -- 8742
,( 7, E,0,0,((45,45),(34,34),( 5, 5),(18,19),(18,18),(14,17)), 1,  9) -- 8743
,( 7, E,0,0,((47,47),(36,36),( 7, 7),(20,21),(20,20),(16,19)), 1,  9) -- 8744
,( 7, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(11,11),( 4, 4)), 1,  9) -- 8745
,( 7, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(13,13),( 6, 6)), 1,  9) -- 8746
,( 7, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(15,15),( 8, 8)), 1,  9) -- 8747
,( 7, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(17,17),(10,10)), 1,  9) -- 8748
,( 7, E,0,0,((44,47),(30,33),( 0, 0),(10,13),( 8,11),( 4, 7)), 1,  8) -- 8749
,( 7, E,0,0,((46,49),(32,35),( 2, 2),(12,15),(10,13),( 6, 9)), 1,  8) -- 8750
,( 7, E,0,0,((48,51),(34,37),( 4, 4),(14,17),(12,15),( 8,11)), 1,  8) -- 8751
,( 7, E,0,0,((50,53),(36,39),( 6, 6),(16,19),(14,17),(10,13)), 1,  8) -- 8752
,( 7, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 8753
,( 7, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 8754
,( 7, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 8755
,( 7, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 8756
,( 7, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(10,13),(99,99)), 1,  8) -- 8757
,( 7, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(12,15),(99,99)), 1,  8) -- 8758
,( 7, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(14,17),(99,99)), 1,  8) -- 8759
,( 7, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(16,19),(99,99)), 1,  8) -- 8760
,( 7, E,0,0,((40,43),(28,31),( 0, 1),(12,15),(14,17),(99,99)), 1,  8) -- 8761
,( 7, E,0,0,((42,45),(30,33),( 2, 3),(14,17),(16,19),(99,99)), 1,  8) -- 8762
,( 7, E,0,0,((44,47),(32,35),( 4, 5),(16,19),(18,21),(99,99)), 1,  8) -- 8763
,( 7, E,0,0,((46,49),(34,37),( 6, 7),(18,21),(20,23),(99,99)), 1,  8) -- 8764
,( 7, E,0,0,((42,45),(28,31),( 0, 1),(14,15),(18,21),(99,99)), 1,  8) -- 8765
,( 7, E,0,0,((44,47),(30,33),( 2, 3),(16,17),(20,23),(99,99)), 1,  8) -- 8766
,( 7, E,0,0,((46,49),(32,35),( 4, 5),(18,19),(22,25),(99,99)), 1,  8) -- 8767
,( 7, E,0,0,((48,51),(34,37),( 6, 7),(20,21),(24,27),(99,99)), 1,  8) -- 8768
,( 7, E,0,0,((48,51),(32,35),( 0, 1),(12,15),(12,15),(99,99)), 1,  7) -- 8769
,( 7, E,0,0,((50,53),(34,37),( 2, 3),(14,17),(14,17),(99,99)), 1,  7) -- 8770
,( 7, E,0,0,((52,55),(36,39),( 4, 5),(16,19),(16,19),(99,99)), 1,  7) -- 8771
,( 7, E,0,0,((54,57),(38,41),( 6, 7),(18,21),(18,21),(99,99)), 1,  7) -- 8772
,( 7, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(16,19),(99,99)), 1,  7) -- 8773
,( 7, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(18,21),(99,99)), 1,  7) -- 8774
,( 7, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(20,23),(99,99)), 1,  7) -- 8775
,( 7, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(22,25),(99,99)), 1,  7) -- 8776
,( 7, E,0,0,((48,51),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 8777
,( 7, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 8778
,( 7, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 8779
,( 7, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 8780
,( 7, E,0,1,((48,51),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 8781
,( 7, E,0,1,((50,53),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 8782
,( 7, E,0,1,((52,55),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 8783
,( 7, E,0,1,((54,57),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 8784
,( 7, E,0,1,((52,55),(34,37),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 8785
,( 7, E,0,1,((54,57),(36,39),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 8786
,( 7, E,0,1,((56,59),(38,41),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 8787
,( 7, E,0,1,((58,61),(40,43),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 8788
,( 7, E,0,1,((48,51),(32,35),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 8789
,( 7, E,0,1,((50,53),(34,37),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 8790
,( 7, E,0,1,((52,55),(36,39),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 8791
,( 7, E,0,1,((54,57),(38,41),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 8792
,( 7, E,0,1,((44,47),(30,33),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 8793
,( 7, E,0,1,((46,49),(32,35),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 8794
,( 7, E,0,1,((48,51),(34,37),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 8795
,( 7, E,0,1,((50,53),(36,39),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 8796
,( 7, E,0,1,((42,45),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 8797
,( 7, E,0,1,((44,47),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 8798
,( 7, E,0,1,((46,49),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 8799
,( 7, E,0,1,((48,51),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 8800
,( 7, E,0,1,((48,51),(30,33),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 8801
,( 7, E,0,1,((50,53),(32,35),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 8802
,( 7, E,0,1,((52,55),(34,37),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 8803
,( 7, E,0,1,((54,57),(36,39),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 8804
,( 7, E,0,1,((40,43),(26,29),( 0, 1),(18,21),(99,99),(99,99)), 1,  5) -- 8805
,( 7, E,0,1,((42,45),(28,31),( 2, 3),(20,23),(99,99),(99,99)), 1,  5) -- 8806
,( 7, E,0,1,((44,47),(30,33),( 4, 5),(22,25),(99,99),(99,99)), 1,  5) -- 8807
,( 7, E,0,1,((46,49),(32,35),( 6, 7),(24,27),(99,99),(99,99)), 1,  5) -- 8808
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 8809
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 8810
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 8811
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 8812
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 8813
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 8814
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 8815
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 8816
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 8817
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 8818
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 8819
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 8820
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 8821
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 8822
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 8823
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 8824
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 8825
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 8826
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 8827
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 8828
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 8829
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 8830
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 8831
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 8832
,( 7, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 8833
,( 7, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 8834
,( 7, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 8835
,( 7, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 8836
,( 7, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 8837
,( 7, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 8838
,( 7, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 8839
,( 7, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 8840
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 8841
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 8842
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 8843
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 8844
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 8845
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 8846
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 8847
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 8848
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 8849
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 8850
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 8851
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 8852
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 8853
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 8854
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 8855
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 8856
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 8857
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 8858
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 8859
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 8860
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 8861
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 8862
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 8863
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 8864
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(17,17),( 8, 8)), 0, 29) -- 8865
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(18,18),( 9, 9)), 0, 29) -- 8866
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(19,19),(10,10)), 0, 29) -- 8867
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(20,20),(11,11)), 0, 29) -- 8868
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(21,21),(12,12)), 0, 29) -- 8869
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(22,22),(13,13)), 0, 29) -- 8870
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(23,23),(14,14)), 0, 29) -- 8871
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(24,24),(15,15)), 0, 29) -- 8872
,( 7, E,0,0,((31,31),(25,25),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 28) -- 8873
,( 7, E,0,0,((32,32),(26,26),( 1, 1),(17,17),(18,18),(10,10)), 0, 28) -- 8874
,( 7, E,0,0,((33,33),(27,27),( 2, 2),(18,18),(19,19),(11,11)), 0, 28) -- 8875
,( 7, E,0,0,((34,34),(28,28),( 3, 3),(19,19),(20,20),(12,12)), 0, 28) -- 8876
,( 7, E,0,0,((35,35),(29,29),( 4, 4),(20,20),(21,21),(13,13)), 0, 28) -- 8877
,( 7, E,0,0,((36,36),(30,30),( 5, 5),(21,21),(22,22),(14,14)), 0, 28) -- 8878
,( 7, E,0,0,((37,37),(31,31),( 6, 6),(22,22),(23,23),(15,15)), 0, 28) -- 8879
,( 7, E,0,0,((38,38),(32,32),( 7, 7),(23,23),(24,24),(16,16)), 0, 28) -- 8880
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 26) -- 8881
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 26) -- 8882
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 26) -- 8883
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 26) -- 8884
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 26) -- 8885
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 26) -- 8886
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 26) -- 8887
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 26) -- 8888
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(15,15),(17,17),( 8, 8)), 0, 25) -- 8889
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(16,16),(18,18),( 9, 9)), 0, 25) -- 8890
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(17,17),(19,19),(10,10)), 0, 25) -- 8891
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(18,18),(20,20),(11,11)), 0, 25) -- 8892
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(19,19),(21,21),(12,12)), 0, 25) -- 8893
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(20,20),(22,22),(13,13)), 0, 25) -- 8894
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(21,21),(23,23),(14,14)), 0, 25) -- 8895
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(22,22),(24,24),(15,15)), 0, 25) -- 8896
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(15,15),(17,17),( 9, 9)), 0, 25) -- 8897
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(16,16),(18,18),(10,10)), 0, 25) -- 8898
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(17,17),(19,19),(11,11)), 0, 25) -- 8899
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(18,18),(20,20),(12,12)), 0, 25) -- 8900
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(19,19),(21,21),(13,13)), 0, 25) -- 8901
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(20,20),(22,22),(14,14)), 0, 25) -- 8902
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(21,21),(23,23),(15,15)), 0, 25) -- 8903
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(22,22),(24,24),(16,16)), 0, 25) -- 8904
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 25) -- 8905
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 25) -- 8906
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 25) -- 8907
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 25) -- 8908
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 25) -- 8909
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 25) -- 8910
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 25) -- 8911
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 25) -- 8912
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 24) -- 8913
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 24) -- 8914
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 24) -- 8915
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 24) -- 8916
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 24) -- 8917
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 24) -- 8918
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 24) -- 8919
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 24) -- 8920
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 24) -- 8921
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(10,10)), 0, 24) -- 8922
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(11,11)), 0, 24) -- 8923
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(12,12)), 0, 24) -- 8924
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(13,13)), 0, 24) -- 8925
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(14,14)), 0, 24) -- 8926
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(15,15)), 0, 24) -- 8927
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(16,16)), 0, 24) -- 8928
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 23) -- 8929
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 23) -- 8930
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 23) -- 8931
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 23) -- 8932
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 23) -- 8933
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 23) -- 8934
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 23) -- 8935
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 23) -- 8936
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(17,17),( 8, 8)), 0, 23) -- 8937
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(18,18),( 9, 9)), 0, 23) -- 8938
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(19,19),(10,10)), 0, 23) -- 8939
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(20,20),(11,11)), 0, 23) -- 8940
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(21,21),(12,12)), 0, 23) -- 8941
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(22,22),(13,13)), 0, 23) -- 8942
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(23,23),(14,14)), 0, 23) -- 8943
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(24,24),(15,15)), 0, 23) -- 8944
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 23) -- 8945
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 23) -- 8946
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 23) -- 8947
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 23) -- 8948
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 23) -- 8949
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 23) -- 8950
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 23) -- 8951
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 23) -- 8952
,( 7, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 22) -- 8953
,( 7, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 22) -- 8954
,( 7, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 22) -- 8955
,( 7, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 22) -- 8956
,( 7, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 22) -- 8957
,( 7, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 22) -- 8958
,( 7, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 22) -- 8959
,( 7, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 22) -- 8960
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 21) -- 8961
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(10,10)), 0, 21) -- 8962
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(11,11)), 0, 21) -- 8963
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(12,12)), 0, 21) -- 8964
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(13,13)), 0, 21) -- 8965
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(14,14)), 0, 21) -- 8966
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(15,15)), 0, 21) -- 8967
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(16,16)), 0, 21) -- 8968
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 8969
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 8970
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 8971
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 8972
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 8973
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 8974
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 8975
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 8976
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 21) -- 8977
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 21) -- 8978
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 21) -- 8979
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 21) -- 8980
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 21) -- 8981
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 21) -- 8982
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 21) -- 8983
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 21) -- 8984
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 8985
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 8986
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 8987
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 8988
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 8989
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 8990
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 8991
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 8992
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 8993
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 8994
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 8995
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 8996
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 8997
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 8998
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 8999
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 9000
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 9001
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 9002
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 9003
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 9004
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 9005
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 9006
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 9007
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 9008
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 19) -- 9009
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 19) -- 9010
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 19) -- 9011
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 19) -- 9012
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 19) -- 9013
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 19) -- 9014
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 19) -- 9015
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 19) -- 9016
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 19) -- 9017
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 19) -- 9018
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 19) -- 9019
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 19) -- 9020
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 19) -- 9021
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 19) -- 9022
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 19) -- 9023
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 19) -- 9024
,( 7, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 9025
,( 7, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 9026
,( 7, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 9027
,( 7, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 9028
,( 7, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 9029
,( 7, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 9030
,( 7, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 9031
,( 7, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 9032
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 19) -- 9033
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 19) -- 9034
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 19) -- 9035
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 19) -- 9036
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 19) -- 9037
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 19) -- 9038
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 19) -- 9039
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 19) -- 9040
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 18) -- 9041
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 18) -- 9042
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 18) -- 9043
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 18) -- 9044
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 18) -- 9045
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 18) -- 9046
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 18) -- 9047
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 18) -- 9048
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 9049
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 9050
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 9051
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 9052
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 9053
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 9054
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 9055
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 9056
,( 7, E,0,0,((30,30),(24,24),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 9057
,( 7, E,0,0,((31,31),(25,25),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 9058
,( 7, E,0,0,((32,32),(26,26),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 9059
,( 7, E,0,0,((33,33),(27,27),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 9060
,( 7, E,0,0,((34,34),(28,28),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 9061
,( 7, E,0,0,((35,35),(29,29),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 9062
,( 7, E,0,0,((36,36),(30,30),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 9063
,( 7, E,0,0,((37,37),(31,31),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 9064
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 18) -- 9065
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 18) -- 9066
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 18) -- 9067
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 18) -- 9068
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 18) -- 9069
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 18) -- 9070
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 18) -- 9071
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 18) -- 9072
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 18) -- 9073
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 18) -- 9074
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 18) -- 9075
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 18) -- 9076
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 18) -- 9077
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 18) -- 9078
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 18) -- 9079
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 18) -- 9080
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 9081
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 9082
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 9083
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 9084
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 9085
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 9086
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 9087
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 9088
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 9089
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 9090
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 9091
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 9092
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 9093
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 9094
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 9095
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 9096
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 17) -- 9097
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 17) -- 9098
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 17) -- 9099
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 17) -- 9100
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 17) -- 9101
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 17) -- 9102
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 17) -- 9103
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 17) -- 9104
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(10,10)), 0, 17) -- 9105
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(11,11)), 0, 17) -- 9106
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(12,12)), 0, 17) -- 9107
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(13,13)), 0, 17) -- 9108
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(14,14)), 0, 17) -- 9109
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(15,15)), 0, 17) -- 9110
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(16,16)), 0, 17) -- 9111
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(17,17)), 0, 17) -- 9112
,( 7, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 9113
,( 7, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 9114
,( 7, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 9115
,( 7, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 9116
,( 7, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 9117
,( 7, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 9118
,( 7, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 9119
,( 7, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 9120
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 16) -- 9121
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 16) -- 9122
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 16) -- 9123
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 16) -- 9124
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 16) -- 9125
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 16) -- 9126
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 16) -- 9127
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 16) -- 9128
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 9129
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 9130
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 9131
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 9132
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 9133
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 9134
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 9135
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 9136
,( 7, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 9137
,( 7, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 9138
,( 7, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 9139
,( 7, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 9140
,( 7, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 9141
,( 7, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 9142
,( 7, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 9143
,( 7, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 9144
,( 7, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 9145
,( 7, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 9146
,( 7, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 9147
,( 7, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 9148
,( 7, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 9149
,( 7, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 9150
,( 7, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 9151
,( 7, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 9152
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(19,19),(11,11)), 0, 16) -- 9153
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(20,20),(12,12)), 0, 16) -- 9154
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(21,21),(13,13)), 0, 16) -- 9155
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(22,22),(14,14)), 0, 16) -- 9156
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(23,23),(15,15)), 0, 16) -- 9157
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(24,24),(16,16)), 0, 16) -- 9158
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(25,25),(17,17)), 0, 16) -- 9159
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(26,26),(18,18)), 0, 16) -- 9160
,( 7, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(19,19),(11,11)), 0, 15) -- 9161
,( 7, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(20,20),(12,12)), 0, 15) -- 9162
,( 7, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(21,21),(13,13)), 0, 15) -- 9163
,( 7, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(22,22),(14,14)), 0, 15) -- 9164
,( 7, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(23,23),(15,15)), 0, 15) -- 9165
,( 7, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(24,24),(16,16)), 0, 15) -- 9166
,( 7, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(25,25),(17,17)), 0, 15) -- 9167
,( 7, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(26,26),(18,18)), 0, 15) -- 9168
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 9169
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 9170
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 9171
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 9172
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 9173
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 9174
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 9175
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 9176
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 15) -- 9177
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 15) -- 9178
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 15) -- 9179
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 15) -- 9180
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 15) -- 9181
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 15) -- 9182
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 15) -- 9183
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 15) -- 9184
,( 7, E,0,0,((28,28),(23,23),( 0, 0),(17,17),(19,19),(10,10)), 0, 15) -- 9185
,( 7, E,0,0,((29,29),(24,24),( 1, 1),(18,18),(20,20),(11,11)), 0, 15) -- 9186
,( 7, E,0,0,((30,30),(25,25),( 2, 2),(19,19),(21,21),(12,12)), 0, 15) -- 9187
,( 7, E,0,0,((31,31),(26,26),( 3, 3),(20,20),(22,22),(13,13)), 0, 15) -- 9188
,( 7, E,0,0,((32,32),(27,27),( 4, 4),(21,21),(23,23),(14,14)), 0, 15) -- 9189
,( 7, E,0,0,((33,33),(28,28),( 5, 5),(22,22),(24,24),(15,15)), 0, 15) -- 9190
,( 7, E,0,0,((34,34),(29,29),( 6, 6),(23,23),(25,25),(16,16)), 0, 15) -- 9191
,( 7, E,0,0,((35,35),(30,30),( 7, 7),(24,24),(26,26),(17,17)), 0, 15) -- 9192
,( 7, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 9193
,( 7, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 9194
,( 7, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 9195
,( 7, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 9196
,( 7, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 9197
,( 7, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 9198
,( 7, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 9199
,( 7, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 9200
,( 7, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 9201
,( 7, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 9202
,( 7, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 9203
,( 7, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 9204
,( 7, E,0,0,((26,29),(22,23),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 9205
,( 7, E,0,0,((28,31),(24,25),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 9206
,( 7, E,0,0,((30,33),(26,27),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 9207
,( 7, E,0,0,((32,35),(28,29),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 9208
,( 7, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(20,20),(10,13)), 0, 14) -- 9209
,( 7, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(22,22),(12,15)), 0, 14) -- 9210
,( 7, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(24,24),(14,17)), 0, 14) -- 9211
,( 7, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(26,26),(16,19)), 0, 14) -- 9212
,( 7, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(10,13)), 0, 13) -- 9213
,( 7, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(12,15)), 0, 13) -- 9214
,( 7, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(14,17)), 0, 13) -- 9215
,( 7, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(16,19)), 0, 13) -- 9216
,( 7, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),( 8, 9)), 0, 13) -- 9217
,( 7, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(10,11)), 0, 13) -- 9218
,( 7, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(12,13)), 0, 13) -- 9219
,( 7, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(14,15)), 0, 13) -- 9220
,( 7, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(10,13)), 0, 12) -- 9221
,( 7, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(12,15)), 0, 12) -- 9222
,( 7, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(14,17)), 0, 12) -- 9223
,( 7, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(16,19)), 0, 12) -- 9224
,( 7, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(22,23),(14,17)), 0, 12) -- 9225
,( 7, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(24,25),(16,19)), 0, 12) -- 9226
,( 7, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(26,27),(18,21)), 0, 12) -- 9227
,( 7, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(28,29),(20,23)), 0, 12) -- 9228
,( 7, E,0,0,((24,27),(20,21),( 0, 1),(18,18),(20,21),(12,15)), 0, 12) -- 9229
,( 7, E,0,0,((26,29),(22,23),( 2, 3),(20,20),(22,23),(14,17)), 0, 12) -- 9230
,( 7, E,0,0,((28,31),(24,25),( 4, 5),(22,22),(24,25),(16,19)), 0, 12) -- 9231
,( 7, E,0,0,((30,33),(26,27),( 6, 7),(24,24),(26,27),(18,21)), 0, 12) -- 9232
,( 7, E,0,0,((24,27),(20,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 12) -- 9233
,( 7, E,0,0,((26,29),(22,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 12) -- 9234
,( 7, E,0,0,((28,31),(24,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 12) -- 9235
,( 7, E,0,0,((30,33),(26,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 12) -- 9236
,( 7, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(12,15)), 0, 11) -- 9237
,( 7, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(14,17)), 0, 11) -- 9238
,( 7, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(16,19)), 0, 11) -- 9239
,( 7, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(18,21)), 0, 11) -- 9240
,( 7, E,0,0,((24,27),(22,23),( 1, 1),(18,19),(22,23),(12,15)), 0, 11) -- 9241
,( 7, E,0,0,((26,29),(24,25),( 3, 3),(20,21),(24,25),(14,17)), 0, 11) -- 9242
,( 7, E,0,0,((28,31),(26,27),( 5, 5),(22,23),(26,27),(16,19)), 0, 11) -- 9243
,( 7, E,0,0,((30,33),(28,29),( 7, 7),(24,25),(28,29),(18,21)), 0, 11) -- 9244
,( 7, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),(10,13)), 0, 11) -- 9245
,( 7, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),(12,15)), 0, 11) -- 9246
,( 7, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(14,17)), 0, 11) -- 9247
,( 7, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(16,19)), 0, 11) -- 9248
,( 7, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(16,19)), 0, 11) -- 9249
,( 7, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(18,21)), 0, 11) -- 9250
,( 7, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(20,23)), 0, 11) -- 9251
,( 7, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(22,23)), 0, 11) -- 9252
,( 7, E,0,0,((25,25),(22,22),( 0, 1),(18,19),(20,21),(10,13)), 0, 11) -- 9253
,( 7, E,0,0,((27,27),(24,24),( 2, 3),(20,21),(22,23),(12,15)), 0, 11) -- 9254
,( 7, E,0,0,((29,29),(26,26),( 4, 5),(22,23),(24,25),(14,17)), 0, 11) -- 9255
,( 7, E,0,0,((31,31),(28,28),( 6, 7),(24,25),(26,27),(16,19)), 0, 11) -- 9256
,( 7, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 9257
,( 7, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 9258
,( 7, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 9259
,( 7, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 9260
,( 7, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),( 8,11)), 0, 10) -- 9261
,( 7, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(10,13)), 0, 10) -- 9262
,( 7, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(12,15)), 0, 10) -- 9263
,( 7, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(14,17)), 0, 10) -- 9264
,( 7, E,0,0,((20,23),(19,19),( 0, 0),(18,19),(22,23),(12,15)), 0, 10) -- 9265
,( 7, E,0,0,((22,25),(21,21),( 2, 2),(20,21),(24,25),(14,17)), 0, 10) -- 9266
,( 7, E,0,0,((24,27),(23,23),( 4, 4),(22,23),(26,27),(16,19)), 0, 10) -- 9267
,( 7, E,0,0,((26,29),(25,25),( 6, 6),(24,25),(28,29),(18,21)), 0, 10) -- 9268
,( 7, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(24,25),(14,17)), 0, 10) -- 9269
,( 7, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(26,27),(16,19)), 0, 10) -- 9270
,( 7, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(28,29),(18,21)), 0, 10) -- 9271
,( 7, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(30,31),(20,23)), 0, 10) -- 9272
,( 7, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(23,23),(12,15)), 0, 10) -- 9273
,( 7, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(25,25),(14,17)), 0, 10) -- 9274
,( 7, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(27,27),(16,19)), 0, 10) -- 9275
,( 7, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(29,29),(18,21)), 0, 10) -- 9276
,( 7, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(18,19),( 6, 9)), 0, 10) -- 9277
,( 7, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(20,21),( 8,11)), 0, 10) -- 9278
,( 7, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(22,23),(10,13)), 0, 10) -- 9279
,( 7, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(24,25),(12,15)), 0, 10) -- 9280
,( 7, E,0,0,((24,27),(22,23),( 0, 1),(18,19),(20,21),( 8, 9)), 0, 10) -- 9281
,( 7, E,0,0,((26,29),(24,25),( 2, 3),(20,21),(22,23),(10,11)), 0, 10) -- 9282
,( 7, E,0,0,((28,31),(26,27),( 4, 5),(22,23),(24,25),(12,13)), 0, 10) -- 9283
,( 7, E,0,0,((30,33),(28,29),( 6, 7),(24,25),(26,27),(14,15)), 0, 10) -- 9284
,( 7, E,0,0,((24,25),(20,21),( 0, 1),(19,19),(24,24),(14,17)), 0, 10) -- 9285
,( 7, E,0,0,((26,27),(22,23),( 2, 3),(21,21),(26,26),(16,19)), 0, 10) -- 9286
,( 7, E,0,0,((28,29),(24,25),( 4, 5),(23,23),(28,28),(18,21)), 0, 10) -- 9287
,( 7, E,0,0,((30,31),(26,27),( 6, 7),(25,25),(30,30),(20,23)), 0, 10) -- 9288
,( 7, E,0,0,((22,22),(19,19),( 0, 0),(18,19),(22,23),(16,19)), 0, 10) -- 9289
,( 7, E,0,0,((24,24),(21,21),( 2, 2),(20,21),(24,25),(18,21)), 0, 10) -- 9290
,( 7, E,0,0,((26,26),(23,23),( 4, 4),(22,23),(26,27),(20,23)), 0, 10) -- 9291
,( 7, E,0,0,((28,28),(25,25),( 6, 6),(24,25),(28,29),(22,23)), 0, 10) -- 9292
,( 7, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 8,11)), 0,  9) -- 9293
,( 7, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),(10,13)), 0,  9) -- 9294
,( 7, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(12,15)), 0,  9) -- 9295
,( 7, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(14,17)), 0,  9) -- 9296
,( 7, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(10,13)), 0,  9) -- 9297
,( 7, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(12,15)), 0,  9) -- 9298
,( 7, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(14,17)), 0,  9) -- 9299
,( 7, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(16,19)), 0,  9) -- 9300
,( 7, E,0,0,((21,21),(18,19),( 0, 1),(20,21),(24,25),(12,15)), 0,  9) -- 9301
,( 7, E,0,0,((23,23),(20,21),( 2, 3),(22,23),(26,27),(14,17)), 0,  9) -- 9302
,( 7, E,0,0,((25,25),(22,23),( 4, 5),(24,25),(28,29),(16,19)), 0,  9) -- 9303
,( 7, E,0,0,((27,27),(24,25),( 6, 7),(26,27),(30,31),(18,21)), 0,  9) -- 9304
,( 7, E,0,0,((20,21),(18,19),( 0, 1),(18,19),(24,25),(12,15)), 0,  9) -- 9305
,( 7, E,0,0,((22,23),(20,21),( 2, 3),(20,21),(26,27),(14,17)), 0,  9) -- 9306
,( 7, E,0,0,((24,25),(22,23),( 4, 5),(22,23),(28,29),(16,19)), 0,  9) -- 9307
,( 7, E,0,0,((26,27),(24,25),( 6, 7),(24,25),(30,31),(18,21)), 0,  9) -- 9308
,( 7, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 9309
,( 7, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 9310
,( 7, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 9311
,( 7, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 9312
,( 7, E,0,0,((20,21),(18,19),( 0, 1),(18,19),(22,23),( 6, 9)), 0,  9) -- 9313
,( 7, E,0,0,((22,23),(20,21),( 2, 3),(20,21),(24,25),( 8,11)), 0,  9) -- 9314
,( 7, E,0,0,((24,25),(22,23),( 4, 5),(22,23),(26,27),(10,13)), 0,  9) -- 9315
,( 7, E,0,0,((26,27),(24,25),( 6, 7),(24,25),(28,29),(12,15)), 0,  9) -- 9316
,( 7, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(20,21),( 4, 7)), 0,  9) -- 9317
,( 7, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(22,23),( 6, 9)), 0,  9) -- 9318
,( 7, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(24,25),( 8,11)), 0,  9) -- 9319
,( 7, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(26,27),(10,13)), 0,  9) -- 9320
,( 7, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 9321
,( 7, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 9322
,( 7, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 9323
,( 7, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 9324
,( 7, E,0,0,((20,23),(20,21),( 0, 1),(18,19),(20,21),( 4, 5)), 0,  9) -- 9325
,( 7, E,0,0,((22,25),(22,23),( 2, 3),(20,21),(22,23),( 6, 7)), 0,  9) -- 9326
,( 7, E,0,0,((24,27),(24,25),( 4, 5),(22,23),(24,25),( 8, 9)), 0,  9) -- 9327
,( 7, E,0,0,((26,29),(26,27),( 6, 7),(24,25),(26,27),(10,11)), 0,  9) -- 9328
,( 7, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(18,19),( 2, 5)), 0,  9) -- 9329
,( 7, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(20,21),( 4, 7)), 0,  9) -- 9330
,( 7, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(22,23),( 6, 9)), 0,  9) -- 9331
,( 7, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(24,25),( 8,11)), 0,  9) -- 9332
,( 7, E,0,0,((23,23),(20,21),( 1, 1),(20,20),(24,24),(10,13)), 0,  9) -- 9333
,( 7, E,0,0,((25,25),(22,23),( 3, 3),(22,22),(26,26),(12,15)), 0,  9) -- 9334
,( 7, E,0,0,((27,27),(24,25),( 5, 5),(24,24),(28,28),(14,17)), 0,  9) -- 9335
,( 7, E,0,0,((29,29),(26,27),( 7, 7),(26,26),(30,30),(16,19)), 0,  9) -- 9336
,( 7, E,0,0,((21,21),(18,19),( 0, 0),(19,19),(24,24),(16,17)), 0,  9) -- 9337
,( 7, E,0,0,((23,23),(20,21),( 2, 2),(21,21),(26,26),(18,19)), 0,  9) -- 9338
,( 7, E,0,0,((25,25),(22,23),( 4, 4),(23,23),(28,28),(20,21)), 0,  9) -- 9339
,( 7, E,0,0,((27,27),(24,25),( 6, 6),(25,25),(30,30),(22,23)), 0,  9) -- 9340
,( 7, E,0,0,((20,23),(20,21),( 1, 1),(20,20),(22,23),( 4, 7)), 0,  9) -- 9341
,( 7, E,0,0,((22,25),(22,23),( 3, 3),(22,22),(24,25),( 6, 9)), 0,  9) -- 9342
,( 7, E,0,0,((24,27),(24,25),( 5, 5),(24,24),(26,27),( 8,11)), 0,  9) -- 9343
,( 7, E,0,0,((26,29),(26,27),( 7, 7),(26,26),(28,29),(10,13)), 0,  9) -- 9344
,( 7, E,0,0,((99,99),(18,19),( 1, 1),(20,20),(23,23),( 8,11)), 0,  9) -- 9345
,( 7, E,0,0,((99,99),(20,21),( 3, 3),(22,22),(25,25),(10,13)), 0,  9) -- 9346
,( 7, E,0,0,((99,99),(22,23),( 5, 5),(24,24),(27,27),(12,15)), 0,  9) -- 9347
,( 7, E,0,0,((99,99),(24,25),( 7, 7),(26,26),(29,29),(14,17)), 0,  9) -- 9348
,( 7, E,0,0,((99,99),(16,19),( 0, 1),(18,21),(22,25),(12,15)), 0,  8) -- 9349
,( 7, E,0,0,((99,99),(18,21),( 2, 3),(20,23),(24,27),(14,17)), 0,  8) -- 9350
,( 7, E,0,0,((99,99),(20,23),( 4, 5),(22,25),(26,29),(16,19)), 0,  8) -- 9351
,( 7, E,0,0,((99,99),(22,25),( 6, 7),(24,27),(28,31),(18,21)), 0,  8) -- 9352
,( 7, E,0,0,((22,25),(18,21),( 0, 1),(18,21),(18,21),(99,99)), 0,  8) -- 9353
,( 7, E,0,0,((24,27),(20,23),( 2, 3),(20,23),(20,23),(99,99)), 0,  8) -- 9354
,( 7, E,0,0,((26,29),(22,25),( 4, 5),(22,25),(22,25),(99,99)), 0,  8) -- 9355
,( 7, E,0,0,((28,31),(24,27),( 6, 7),(24,27),(24,27),(99,99)), 0,  8) -- 9356
,( 7, E,0,0,((99,99),(16,19),( 0, 1),(18,21),(26,29),(17,17)), 0,  8) -- 9357
,( 7, E,0,0,((99,99),(18,21),( 2, 3),(20,23),(28,31),(19,19)), 0,  8) -- 9358
,( 7, E,0,0,((99,99),(20,23),( 4, 5),(22,25),(30,33),(21,21)), 0,  8) -- 9359
,( 7, E,0,0,((99,99),(22,25),( 6, 7),(24,27),(32,35),(23,23)), 0,  8) -- 9360
,( 7, E,0,0,((99,99),(16,17),( 0, 1),(18,21),(18,21),(99,99)), 0,  7) -- 9361
,( 7, E,0,0,((99,99),(18,19),( 2, 3),(20,23),(20,23),(99,99)), 0,  7) -- 9362
,( 7, E,0,0,((99,99),(20,21),( 4, 5),(22,25),(22,25),(99,99)), 0,  7) -- 9363
,( 7, E,0,0,((99,99),(22,23),( 6, 7),(24,27),(24,27),(99,99)), 0,  7) -- 9364
,( 7, E,0,1,((99,99),(16,19),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 9365
,( 7, E,0,1,((99,99),(18,21),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 9366
,( 7, E,0,1,((99,99),(20,23),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 9367
,( 7, E,0,1,((99,99),(22,25),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 9368
,( 7, E,0,1,((99,99),(18,21),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 9369
,( 7, E,0,1,((99,99),(20,23),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 9370
,( 7, E,0,1,((99,99),(22,25),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 9371
,( 7, E,0,1,((99,99),(24,27),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 9372
,( 7, E,0,1,((22,25),(20,23),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 9373
,( 7, E,0,1,((24,27),(22,25),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 9374
,( 7, E,0,1,((26,29),(24,27),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 9375
,( 7, E,0,1,((28,31),(26,29),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 9376
,( 7, E,0,1,((99,99),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 9377
,( 7, E,0,1,((99,99),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 9378
,( 7, E,0,1,((99,99),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 9379
,( 7, E,0,1,((99,99),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 9380
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 9381
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 9382
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 9383
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 9384
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 9385
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 9386
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 9387
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 9388
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 9389
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 9390
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 9391
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 9392
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 9393
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 9394
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 9395
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 9396
,( 8, E,0,0,((32,32),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 9397
,( 8, E,0,0,((33,33),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 9398
,( 8, E,0,0,((34,34),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 9399
,( 8, E,0,0,((35,35),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 9400
,( 8, E,0,0,((36,36),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 9401
,( 8, E,0,0,((37,37),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 9402
,( 8, E,0,0,((38,38),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 9403
,( 8, E,0,0,((39,39),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 9404
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 9405
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 9406
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 9407
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 9408
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 9409
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 9410
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 9411
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 9412
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 9413
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 9414
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 9415
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 9416
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 9417
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 9418
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 9419
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 9420
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 31) -- 9421
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 1, 31) -- 9422
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 1, 31) -- 9423
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 1, 31) -- 9424
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 1, 31) -- 9425
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 1, 31) -- 9426
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 1, 31) -- 9427
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 1, 31) -- 9428
,( 8, E,0,0,((32,32),(23,23),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 9429
,( 8, E,0,0,((33,33),(24,24),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 9430
,( 8, E,0,0,((34,34),(25,25),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 9431
,( 8, E,0,0,((35,35),(26,26),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 9432
,( 8, E,0,0,((36,36),(27,27),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 9433
,( 8, E,0,0,((37,37),(28,28),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 9434
,( 8, E,0,0,((38,38),(29,29),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 9435
,( 8, E,0,0,((39,39),(30,30),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 9436
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 31) -- 9437
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 31) -- 9438
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 1, 31) -- 9439
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 1, 31) -- 9440
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 1, 31) -- 9441
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 1, 31) -- 9442
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 1, 31) -- 9443
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 1, 31) -- 9444
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 31) -- 9445
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 31) -- 9446
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 31) -- 9447
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 31) -- 9448
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 31) -- 9449
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 31) -- 9450
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 31) -- 9451
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 31) -- 9452
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 30) -- 9453
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 30) -- 9454
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 30) -- 9455
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 30) -- 9456
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 30) -- 9457
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 30) -- 9458
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 30) -- 9459
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 30) -- 9460
,( 8, E,0,0,((32,32),(23,23),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 29) -- 9461
,( 8, E,0,0,((33,33),(24,24),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 29) -- 9462
,( 8, E,0,0,((34,34),(25,25),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 29) -- 9463
,( 8, E,0,0,((35,35),(26,26),( 3, 3),(18,18),(18,18),(10,10)), 1, 29) -- 9464
,( 8, E,0,0,((36,36),(27,27),( 4, 4),(19,19),(19,19),(11,11)), 1, 29) -- 9465
,( 8, E,0,0,((37,37),(28,28),( 5, 5),(20,20),(20,20),(12,12)), 1, 29) -- 9466
,( 8, E,0,0,((38,38),(29,29),( 6, 6),(21,21),(21,21),(13,13)), 1, 29) -- 9467
,( 8, E,0,0,((39,39),(30,30),( 7, 7),(22,22),(22,22),(14,14)), 1, 29) -- 9468
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 28) -- 9469
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 28) -- 9470
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 28) -- 9471
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 28) -- 9472
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 28) -- 9473
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 28) -- 9474
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 28) -- 9475
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 28) -- 9476
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 26) -- 9477
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 26) -- 9478
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 26) -- 9479
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 26) -- 9480
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 26) -- 9481
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 26) -- 9482
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 26) -- 9483
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 26) -- 9484
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 24) -- 9485
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 24) -- 9486
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 24) -- 9487
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 24) -- 9488
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 24) -- 9489
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 24) -- 9490
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 24) -- 9491
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 24) -- 9492
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 23) -- 9493
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 23) -- 9494
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 23) -- 9495
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 23) -- 9496
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 23) -- 9497
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 23) -- 9498
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 23) -- 9499
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 23) -- 9500
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 9501
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 9502
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 9503
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 9504
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 9505
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 9506
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 9507
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 9508
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 22) -- 9509
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 22) -- 9510
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 22) -- 9511
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 22) -- 9512
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 22) -- 9513
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 22) -- 9514
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 22) -- 9515
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 22) -- 9516
,( 8, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 22) -- 9517
,( 8, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 22) -- 9518
,( 8, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 22) -- 9519
,( 8, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 22) -- 9520
,( 8, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 22) -- 9521
,( 8, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 22) -- 9522
,( 8, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 22) -- 9523
,( 8, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 22) -- 9524
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 22) -- 9525
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 22) -- 9526
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 22) -- 9527
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 22) -- 9528
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 22) -- 9529
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 22) -- 9530
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 22) -- 9531
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 22) -- 9532
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 21) -- 9533
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 21) -- 9534
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 21) -- 9535
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 21) -- 9536
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 21) -- 9537
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 21) -- 9538
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 21) -- 9539
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 21) -- 9540
,( 8, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 9541
,( 8, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 9542
,( 8, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 9543
,( 8, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 9544
,( 8, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 9545
,( 8, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 9546
,( 8, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 9547
,( 8, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 9548
,( 8, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 20) -- 9549
,( 8, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 20) -- 9550
,( 8, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 20) -- 9551
,( 8, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 20) -- 9552
,( 8, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 20) -- 9553
,( 8, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 20) -- 9554
,( 8, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 20) -- 9555
,( 8, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 20) -- 9556
,( 8, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 20) -- 9557
,( 8, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 20) -- 9558
,( 8, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 20) -- 9559
,( 8, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 20) -- 9560
,( 8, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 20) -- 9561
,( 8, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 20) -- 9562
,( 8, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 20) -- 9563
,( 8, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 20) -- 9564
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 9565
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 9566
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 9567
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 9568
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 9569
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 9570
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 9571
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 9572
,( 8, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 19) -- 9573
,( 8, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 19) -- 9574
,( 8, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 19) -- 9575
,( 8, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 19) -- 9576
,( 8, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 19) -- 9577
,( 8, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 19) -- 9578
,( 8, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 19) -- 9579
,( 8, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 19) -- 9580
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 9581
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 9582
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 9583
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 9584
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 9585
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 9586
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 9587
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 9588
,( 8, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 9589
,( 8, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 9590
,( 8, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 9591
,( 8, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 9592
,( 8, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 9593
,( 8, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 9594
,( 8, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 9595
,( 8, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 9596
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 19) -- 9597
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 19) -- 9598
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 19) -- 9599
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 19) -- 9600
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 19) -- 9601
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 19) -- 9602
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 19) -- 9603
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 19) -- 9604
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 9605
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 9606
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 9607
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 9608
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 9609
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 9610
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 9611
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 9612
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 18) -- 9613
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 18) -- 9614
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 18) -- 9615
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 18) -- 9616
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 18) -- 9617
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 18) -- 9618
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 18) -- 9619
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 18) -- 9620
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 9621
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 9622
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 9623
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 9624
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 9625
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 9626
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 9627
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 9628
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 9629
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 9630
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 9631
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 9632
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 9633
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 9634
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 9635
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 9636
,( 8, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 9637
,( 8, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 9638
,( 8, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 9639
,( 8, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 9640
,( 8, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 9641
,( 8, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 9642
,( 8, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 9643
,( 8, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 9644
,( 8, E,0,0,((34,34),(24,24),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 9645
,( 8, E,0,0,((35,35),(25,25),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 9646
,( 8, E,0,0,((36,36),(26,26),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 9647
,( 8, E,0,0,((37,37),(27,27),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 9648
,( 8, E,0,0,((38,38),(28,28),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 9649
,( 8, E,0,0,((39,39),(29,29),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 9650
,( 8, E,0,0,((40,40),(30,30),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 9651
,( 8, E,0,0,((41,41),(31,31),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 9652
,( 8, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 9653
,( 8, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 9654
,( 8, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 9655
,( 8, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 9656
,( 8, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 9657
,( 8, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 9658
,( 8, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 9659
,( 8, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 9660
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 9661
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 9662
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 9663
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 9664
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 9665
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 9666
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 9667
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 9668
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 9669
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 9670
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 9671
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 9672
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 9673
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 9674
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 9675
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 9676
,( 8, E,0,0,((34,34),(24,24),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 9677
,( 8, E,0,0,((35,35),(25,25),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 9678
,( 8, E,0,0,((36,36),(26,26),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 9679
,( 8, E,0,0,((37,37),(27,27),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 9680
,( 8, E,0,0,((38,38),(28,28),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 9681
,( 8, E,0,0,((39,39),(29,29),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 9682
,( 8, E,0,0,((40,40),(30,30),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 9683
,( 8, E,0,0,((41,41),(31,31),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 9684
,( 8, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 9685
,( 8, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 9686
,( 8, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 9687
,( 8, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 9688
,( 8, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 9689
,( 8, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 9690
,( 8, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 9691
,( 8, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 9692
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 9693
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 9694
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 9695
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 9696
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 9697
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 9698
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 9699
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 9700
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 9701
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 9702
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 9703
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 9704
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 9705
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 9706
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 9707
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 9708
,( 8, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 9709
,( 8, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 9710
,( 8, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 9711
,( 8, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 9712
,( 8, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 9713
,( 8, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 9714
,( 8, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 9715
,( 8, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 9716
,( 8, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 16) -- 9717
,( 8, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 16) -- 9718
,( 8, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 16) -- 9719
,( 8, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 16) -- 9720
,( 8, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 16) -- 9721
,( 8, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 16) -- 9722
,( 8, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 16) -- 9723
,( 8, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 16) -- 9724
,( 8, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 16) -- 9725
,( 8, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 16) -- 9726
,( 8, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 16) -- 9727
,( 8, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 16) -- 9728
,( 8, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 16) -- 9729
,( 8, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 16) -- 9730
,( 8, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 16) -- 9731
,( 8, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 16) -- 9732
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 15) -- 9733
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 15) -- 9734
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 15) -- 9735
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 15) -- 9736
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 15) -- 9737
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 15) -- 9738
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 15) -- 9739
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 15) -- 9740
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 9741
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 9742
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 9743
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 9744
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 9745
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 9746
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 9747
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 9748
,( 8, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 15) -- 9749
,( 8, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 15) -- 9750
,( 8, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 15) -- 9751
,( 8, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 15) -- 9752
,( 8, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 15) -- 9753
,( 8, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 15) -- 9754
,( 8, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 15) -- 9755
,( 8, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 15) -- 9756
,( 8, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 9757
,( 8, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 9758
,( 8, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 9759
,( 8, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 9760
,( 8, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 9761
,( 8, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 9762
,( 8, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 9763
,( 8, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 9764
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 9765
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 9766
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 9767
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 9768
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 9769
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 9770
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 9771
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 9772
,( 8, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 9773
,( 8, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 9774
,( 8, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 9775
,( 8, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 9776
,( 8, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 9777
,( 8, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 9778
,( 8, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 9779
,( 8, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 9780
,( 8, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 9781
,( 8, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 9782
,( 8, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 9783
,( 8, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 9784
,( 8, E,0,0,((36,39),(26,27),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 9785
,( 8, E,0,0,((38,41),(28,29),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 9786
,( 8, E,0,0,((40,43),(30,31),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 9787
,( 8, E,0,0,((42,45),(32,33),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 9788
,( 8, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 13) -- 9789
,( 8, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 13) -- 9790
,( 8, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 13) -- 9791
,( 8, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 13) -- 9792
,( 8, E,0,0,((38,38),(27,27),( 1, 1),(15,15),(14,15),( 4, 7)), 1, 13) -- 9793
,( 8, E,0,0,((40,40),(29,29),( 3, 3),(17,17),(16,17),( 6, 9)), 1, 13) -- 9794
,( 8, E,0,0,((42,42),(31,31),( 5, 5),(19,19),(18,19),( 8,11)), 1, 13) -- 9795
,( 8, E,0,0,((44,44),(33,33),( 7, 7),(21,21),(20,21),(10,13)), 1, 13) -- 9796
,( 8, E,0,0,((38,41),(28,28),( 1, 1),(15,15),(14,15),( 4, 7)), 1, 12) -- 9797
,( 8, E,0,0,((40,43),(30,30),( 3, 3),(17,17),(16,17),( 6, 9)), 1, 12) -- 9798
,( 8, E,0,0,((42,45),(32,32),( 5, 5),(19,19),(18,19),( 8,11)), 1, 12) -- 9799
,( 8, E,0,0,((44,47),(34,34),( 7, 7),(21,21),(20,21),(10,13)), 1, 12) -- 9800
,( 8, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 9801
,( 8, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 9802
,( 8, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 9803
,( 8, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 9804
,( 8, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(13,13),( 6, 6)), 1, 12) -- 9805
,( 8, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(15,15),( 8, 8)), 1, 12) -- 9806
,( 8, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(17,17),(10,10)), 1, 12) -- 9807
,( 8, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(19,19),(12,12)), 1, 12) -- 9808
,( 8, E,0,0,((38,41),(26,27),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 11) -- 9809
,( 8, E,0,0,((40,43),(28,29),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 11) -- 9810
,( 8, E,0,0,((42,45),(30,31),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 11) -- 9811
,( 8, E,0,0,((44,47),(32,33),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 11) -- 9812
,( 8, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 11) -- 9813
,( 8, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 11) -- 9814
,( 8, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 11) -- 9815
,( 8, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(18,18),( 8,11)), 1, 11) -- 9816
,( 8, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 7)), 1, 11) -- 9817
,( 8, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8, 9)), 1, 11) -- 9818
,( 8, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,11)), 1, 11) -- 9819
,( 8, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,13)), 1, 11) -- 9820
,( 8, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 9821
,( 8, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 9822
,( 8, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),(10,13)), 1, 11) -- 9823
,( 8, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(12,15)), 1, 11) -- 9824
,( 8, E,0,0,((38,41),(28,29),( 0, 1),(13,13),(10,11),( 0, 3)), 1, 11) -- 9825
,( 8, E,0,0,((40,43),(30,31),( 2, 3),(15,15),(12,13),( 2, 5)), 1, 11) -- 9826
,( 8, E,0,0,((42,45),(32,33),( 4, 5),(17,17),(14,15),( 4, 7)), 1, 11) -- 9827
,( 8, E,0,0,((44,47),(34,35),( 6, 7),(19,19),(16,17),( 6, 9)), 1, 11) -- 9828
,( 8, E,0,0,((38,41),(28,29),( 1, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 9829
,( 8, E,0,0,((40,43),(30,31),( 3, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 9830
,( 8, E,0,0,((42,45),(32,33),( 5, 5),(18,19),(18,19),(10,13)), 1, 11) -- 9831
,( 8, E,0,0,((44,47),(34,35),( 7, 7),(20,21),(20,21),(12,15)), 1, 11) -- 9832
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(11,11),( 0, 3)), 1, 11) -- 9833
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(13,13),( 2, 5)), 1, 11) -- 9834
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(15,15),( 4, 7)), 1, 11) -- 9835
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(17,17),( 6, 9)), 1, 11) -- 9836
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(10,11),( 2, 5)), 1, 10) -- 9837
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(12,13),( 4, 7)), 1, 10) -- 9838
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(14,15),( 6, 9)), 1, 10) -- 9839
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(16,17),( 8,11)), 1, 10) -- 9840
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(13,13),(12,12),( 4, 7)), 1, 10) -- 9841
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(15,15),(14,14),( 6, 9)), 1, 10) -- 9842
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(17,17),(16,16),( 8,11)), 1, 10) -- 9843
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(19,19),(18,18),(10,13)), 1, 10) -- 9844
,( 8, E,0,0,((42,42),(29,29),( 0, 1),(14,15),(12,13),( 4, 7)), 1, 10) -- 9845
,( 8, E,0,0,((44,44),(31,31),( 2, 3),(16,17),(14,15),( 6, 9)), 1, 10) -- 9846
,( 8, E,0,0,((46,46),(33,33),( 4, 5),(18,19),(16,17),( 8,11)), 1, 10) -- 9847
,( 8, E,0,0,((48,48),(35,35),( 6, 7),(20,21),(18,19),(10,13)), 1, 10) -- 9848
,( 8, E,0,0,((42,43),(30,30),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 10) -- 9849
,( 8, E,0,0,((44,45),(32,32),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 10) -- 9850
,( 8, E,0,0,((46,47),(34,34),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 10) -- 9851
,( 8, E,0,0,((48,49),(36,36),( 7, 7),(20,21),(18,19),( 8,11)), 1, 10) -- 9852
,( 8, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1, 10) -- 9853
,( 8, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1, 10) -- 9854
,( 8, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1, 10) -- 9855
,( 8, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1, 10) -- 9856
,( 8, E,0,0,((38,41),(27,27),( 0, 0),(14,14),(12,13),( 6, 9)), 1, 10) -- 9857
,( 8, E,0,0,((40,43),(29,29),( 2, 2),(16,16),(14,15),( 8,11)), 1, 10) -- 9858
,( 8, E,0,0,((42,45),(31,31),( 4, 4),(18,18),(16,17),(10,13)), 1, 10) -- 9859
,( 8, E,0,0,((44,47),(33,33),( 6, 6),(20,20),(18,19),(12,15)), 1, 10) -- 9860
,( 8, E,0,0,((42,45),(30,30),( 1, 1),(14,14),(10,11),( 0, 3)), 1, 10) -- 9861
,( 8, E,0,0,((44,47),(32,32),( 3, 3),(16,16),(12,13),( 2, 5)), 1, 10) -- 9862
,( 8, E,0,0,((46,49),(34,34),( 5, 5),(18,18),(14,15),( 4, 7)), 1, 10) -- 9863
,( 8, E,0,0,((48,51),(36,36),( 7, 7),(20,20),(16,17),( 6, 9)), 1, 10) -- 9864
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(12,13),( 8, 9)), 1, 10) -- 9865
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(14,15),(10,11)), 1, 10) -- 9866
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(16,17),(12,13)), 1, 10) -- 9867
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(18,19),(14,15)), 1, 10) -- 9868
,( 8, E,0,0,((40,43),(28,29),( 0, 0),(12,13),( 8, 9),( 0, 3)), 1, 10) -- 9869
,( 8, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(10,11),( 2, 5)), 1, 10) -- 9870
,( 8, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(12,13),( 4, 7)), 1, 10) -- 9871
,( 8, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(14,15),( 6, 9)), 1, 10) -- 9872
,( 8, E,0,0,((38,41),(28,29),( 0, 1),(14,14),(11,11),( 2, 5)), 1, 10) -- 9873
,( 8, E,0,0,((40,43),(30,31),( 2, 3),(16,16),(13,13),( 4, 7)), 1, 10) -- 9874
,( 8, E,0,0,((42,45),(32,33),( 4, 5),(18,18),(15,15),( 6, 9)), 1, 10) -- 9875
,( 8, E,0,0,((44,47),(34,35),( 6, 7),(20,20),(17,17),( 8,11)), 1, 10) -- 9876
,( 8, E,0,0,((42,42),(29,29),( 0, 1),(14,15),(12,12),( 2, 3)), 1, 10) -- 9877
,( 8, E,0,0,((44,44),(31,31),( 2, 3),(16,17),(14,14),( 4, 5)), 1, 10) -- 9878
,( 8, E,0,0,((46,46),(33,33),( 4, 5),(18,19),(16,16),( 6, 7)), 1, 10) -- 9879
,( 8, E,0,0,((48,48),(35,35),( 6, 7),(20,21),(18,18),( 8, 9)), 1, 10) -- 9880
,( 8, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),( 6, 9)), 1,  9) -- 9881
,( 8, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),( 8,11)), 1,  9) -- 9882
,( 8, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(10,13)), 1,  9) -- 9883
,( 8, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(12,15)), 1,  9) -- 9884
,( 8, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1,  9) -- 9885
,( 8, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 8,11)), 1,  9) -- 9886
,( 8, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(10,13)), 1,  9) -- 9887
,( 8, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(12,15)), 1,  9) -- 9888
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(12,13),( 8,11)), 1,  9) -- 9889
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(14,15),(10,13)), 1,  9) -- 9890
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(16,17),(12,15)), 1,  9) -- 9891
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(18,19),(14,17)), 1,  9) -- 9892
,( 8, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 9893
,( 8, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 9894
,( 8, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 9895
,( 8, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 9896
,( 8, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 9897
,( 8, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 9898
,( 8, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(10,13)), 1,  9) -- 9899
,( 8, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(12,15)), 1,  9) -- 9900
,( 8, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(11,11),( 4, 7)), 1,  9) -- 9901
,( 8, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(13,13),( 6, 9)), 1,  9) -- 9902
,( 8, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(15,15),( 8,11)), 1,  9) -- 9903
,( 8, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(17,17),(10,13)), 1,  9) -- 9904
,( 8, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 9905
,( 8, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 9906
,( 8, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 9907
,( 8, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 9908
,( 8, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(14,15),( 8,11)), 1,  9) -- 9909
,( 8, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(16,17),(10,13)), 1,  9) -- 9910
,( 8, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(18,19),(12,15)), 1,  9) -- 9911
,( 8, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(20,21),(14,17)), 1,  9) -- 9912
,( 8, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 8,11)), 1,  9) -- 9913
,( 8, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(10,13)), 1,  9) -- 9914
,( 8, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(12,15)), 1,  9) -- 9915
,( 8, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(14,17)), 1,  9) -- 9916
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(12,13),(10,13)), 1,  9) -- 9917
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(14,15),(12,15)), 1,  9) -- 9918
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(16,17),(14,17)), 1,  9) -- 9919
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(18,19),(16,19)), 1,  9) -- 9920
,( 8, E,0,0,((42,43),(29,29),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 9921
,( 8, E,0,0,((44,45),(31,31),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 9922
,( 8, E,0,0,((46,47),(33,33),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 9923
,( 8, E,0,0,((48,49),(35,35),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 9924
,( 8, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),(10,13)), 1,  9) -- 9925
,( 8, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),(12,15)), 1,  9) -- 9926
,( 8, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(14,17)), 1,  9) -- 9927
,( 8, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(16,19)), 1,  9) -- 9928
,( 8, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),(12,15)), 1,  9) -- 9929
,( 8, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),(14,17)), 1,  9) -- 9930
,( 8, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(16,19)), 1,  9) -- 9931
,( 8, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(18,21)), 1,  9) -- 9932
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(10,11),( 0, 1)), 1,  9) -- 9933
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(12,13),( 2, 3)), 1,  9) -- 9934
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(14,15),( 4, 5)), 1,  9) -- 9935
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(16,17),( 6, 7)), 1,  9) -- 9936
,( 8, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(11,11),(10,13)), 1,  9) -- 9937
,( 8, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(13,13),(12,15)), 1,  9) -- 9938
,( 8, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(15,15),(14,17)), 1,  9) -- 9939
,( 8, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(17,17),(16,19)), 1,  9) -- 9940
,( 8, E,0,0,((42,43),(29,29),( 0, 1),(14,14),(10,11),( 2, 5)), 1,  9) -- 9941
,( 8, E,0,0,((44,45),(31,31),( 2, 3),(16,16),(12,13),( 4, 7)), 1,  9) -- 9942
,( 8, E,0,0,((46,47),(33,33),( 4, 5),(18,18),(14,15),( 6, 9)), 1,  9) -- 9943
,( 8, E,0,0,((48,49),(35,35),( 6, 7),(20,20),(16,17),( 8,11)), 1,  9) -- 9944
,( 8, E,0,0,((40,43),(29,29),( 0, 1),(14,15),(14,14),( 8, 9)), 1,  9) -- 9945
,( 8, E,0,0,((42,45),(31,31),( 2, 3),(16,17),(16,16),(10,11)), 1,  9) -- 9946
,( 8, E,0,0,((44,47),(33,33),( 4, 5),(18,19),(18,18),(12,13)), 1,  9) -- 9947
,( 8, E,0,0,((46,49),(35,35),( 6, 7),(20,21),(20,20),(14,15)), 1,  9) -- 9948
,( 8, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(10,13),( 7, 7)), 1,  8) -- 9949
,( 8, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(12,15),( 9, 9)), 1,  8) -- 9950
,( 8, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(14,17),(11,11)), 1,  8) -- 9951
,( 8, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(16,19),(13,13)), 1,  8) -- 9952
,( 8, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(14,17),(13,13)), 1,  8) -- 9953
,( 8, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(16,19),(15,15)), 1,  8) -- 9954
,( 8, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(18,21),(17,17)), 1,  8) -- 9955
,( 8, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(20,23),(19,19)), 1,  8) -- 9956
,( 8, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 6, 9),( 2, 5)), 1,  8) -- 9957
,( 8, E,0,0,((46,49),(32,35),( 2, 3),(12,15),( 8,11),( 4, 7)), 1,  8) -- 9958
,( 8, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(10,13),( 6, 9)), 1,  8) -- 9959
,( 8, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(12,15),( 8,11)), 1,  8) -- 9960
,( 8, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(14,17)), 1,  8) -- 9961
,( 8, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(16,19)), 1,  8) -- 9962
,( 8, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(18,21)), 1,  8) -- 9963
,( 8, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(20,23)), 1,  8) -- 9964
,( 8, E,0,0,((48,49),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  7) -- 9965
,( 8, E,0,0,((50,51),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  7) -- 9966
,( 8, E,0,0,((52,53),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  7) -- 9967
,( 8, E,0,0,((54,55),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  7) -- 9968
,( 8, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(18,19),(99,99)), 1,  7) -- 9969
,( 8, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(20,21),(99,99)), 1,  7) -- 9970
,( 8, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(22,23),(99,99)), 1,  7) -- 9971
,( 8, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(24,25),(99,99)), 1,  7) -- 9972
,( 8, E,0,0,((48,51),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 9973
,( 8, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 9974
,( 8, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 9975
,( 8, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 9976
,( 8, E,0,1,((50,53),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 9977
,( 8, E,0,1,((52,55),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 9978
,( 8, E,0,1,((54,57),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 9979
,( 8, E,0,1,((56,59),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 9980
,( 8, E,0,1,((48,51),(30,33),( 0, 1),(14,17),(99,99),(99,99)), 1,  7) -- 9981
,( 8, E,0,1,((50,53),(32,35),( 2, 3),(16,19),(99,99),(99,99)), 1,  7) -- 9982
,( 8, E,0,1,((52,55),(34,37),( 4, 5),(18,21),(99,99),(99,99)), 1,  7) -- 9983
,( 8, E,0,1,((54,57),(36,39),( 6, 7),(20,23),(99,99),(99,99)), 1,  7) -- 9984
,( 8, E,0,1,((44,47),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 9985
,( 8, E,0,1,((46,49),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 9986
,( 8, E,0,1,((48,51),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 9987
,( 8, E,0,1,((50,53),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 9988
,( 8, E,0,1,((52,55),(32,35),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 9989
,( 8, E,0,1,((54,57),(34,37),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 9990
,( 8, E,0,1,((56,59),(36,39),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 9991
,( 8, E,0,1,((58,61),(38,41),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 9992
,( 8, E,0,1,((48,51),(32,35),( 0, 1),( 8,11),(99,99),(99,99)), 1,  6) -- 9993
,( 8, E,0,1,((50,53),(34,37),( 2, 3),(10,13),(99,99),(99,99)), 1,  6) -- 9994
,( 8, E,0,1,((52,55),(36,39),( 4, 5),(12,15),(99,99),(99,99)), 1,  6) -- 9995
,( 8, E,0,1,((54,57),(38,41),( 6, 7),(14,17),(99,99),(99,99)), 1,  6) -- 9996
,( 8, E,0,1,((38,41),(26,27),( 0, 1),(16,19),(99,99),(99,99)), 1,  5) -- 9997
,( 8, E,0,1,((40,43),(28,29),( 2, 3),(18,21),(99,99),(99,99)), 1,  5) -- 9998
,( 8, E,0,1,((42,45),(30,31),( 4, 5),(20,23),(99,99),(99,99)), 1,  5) -- 9999
,( 8, E,0,1,((44,47),(32,33),( 6, 7),(22,25),(99,99),(99,99)), 1,  5) -- 10000
,( 8, E,0,1,((40,43),(26,29),( 0, 1),(24,25),(99,99),(99,99)), 1,  5) -- 10001
,( 8, E,0,1,((42,45),(28,31),( 2, 3),(26,27),(99,99),(99,99)), 1,  5) -- 10002
,( 8, E,0,1,((44,47),(30,33),( 4, 5),(28,29),(99,99),(99,99)), 1,  5) -- 10003
,( 8, E,0,1,((46,49),(32,35),( 6, 7),(30,31),(99,99),(99,99)), 1,  5) -- 10004
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 10005
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 10006
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 10007
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 10008
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 10009
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 10010
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 10011
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 10012
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 10013
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 10014
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 10015
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 10016
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 10017
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 10018
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 10019
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 10020
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 10021
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 10022
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 10023
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 10024
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 10025
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 10026
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 10027
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 10028
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 10029
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 10030
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 10031
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 10032
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 10033
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 10034
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 10035
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 10036
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 10037
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 10038
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 10039
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 10040
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 10041
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 10042
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 10043
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 10044
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 10045
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 10046
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 10047
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 10048
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 10049
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 10050
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 10051
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 10052
,( 8, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 10053
,( 8, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 10054
,( 8, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 10055
,( 8, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 10056
,( 8, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 10057
,( 8, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 10058
,( 8, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 10059
,( 8, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 10060
,( 8, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 10061
,( 8, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 10062
,( 8, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 10063
,( 8, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 10064
,( 8, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 10065
,( 8, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 10066
,( 8, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 10067
,( 8, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 10068
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 30) -- 10069
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 30) -- 10070
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 30) -- 10071
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 30) -- 10072
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 30) -- 10073
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 30) -- 10074
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 30) -- 10075
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 30) -- 10076
,( 8, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 30) -- 10077
,( 8, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 30) -- 10078
,( 8, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 30) -- 10079
,( 8, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 30) -- 10080
,( 8, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 30) -- 10081
,( 8, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 30) -- 10082
,( 8, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 30) -- 10083
,( 8, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 30) -- 10084
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 27) -- 10085
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 27) -- 10086
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 27) -- 10087
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 27) -- 10088
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 27) -- 10089
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 27) -- 10090
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 27) -- 10091
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 27) -- 10092
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 25) -- 10093
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 25) -- 10094
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 25) -- 10095
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 25) -- 10096
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 25) -- 10097
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 25) -- 10098
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 25) -- 10099
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 25) -- 10100
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 24) -- 10101
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 24) -- 10102
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 24) -- 10103
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 24) -- 10104
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 24) -- 10105
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 24) -- 10106
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 24) -- 10107
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 24) -- 10108
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 24) -- 10109
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 24) -- 10110
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 24) -- 10111
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 24) -- 10112
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 24) -- 10113
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 24) -- 10114
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 24) -- 10115
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 24) -- 10116
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 24) -- 10117
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 24) -- 10118
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 24) -- 10119
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 24) -- 10120
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 24) -- 10121
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 24) -- 10122
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 24) -- 10123
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 24) -- 10124
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 23) -- 10125
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 23) -- 10126
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 23) -- 10127
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 23) -- 10128
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 23) -- 10129
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 23) -- 10130
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 23) -- 10131
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 23) -- 10132
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 23) -- 10133
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 23) -- 10134
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 23) -- 10135
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 23) -- 10136
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 23) -- 10137
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 23) -- 10138
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 23) -- 10139
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 23) -- 10140
,( 8, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 21) -- 10141
,( 8, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 21) -- 10142
,( 8, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 21) -- 10143
,( 8, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 21) -- 10144
,( 8, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 21) -- 10145
,( 8, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 21) -- 10146
,( 8, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 21) -- 10147
,( 8, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 21) -- 10148
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 10149
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 10150
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 10151
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 10152
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 10153
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 10154
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 10155
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 10156
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 10157
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 10158
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 10159
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 10160
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 10161
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 10162
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 10163
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 10164
,( 8, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 10165
,( 8, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 10166
,( 8, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 10167
,( 8, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 10168
,( 8, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 10169
,( 8, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 10170
,( 8, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 10171
,( 8, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 10172
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 20) -- 10173
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 20) -- 10174
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 20) -- 10175
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 20) -- 10176
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 20) -- 10177
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 20) -- 10178
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 20) -- 10179
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 20) -- 10180
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 10181
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 10182
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 10183
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 10184
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 10185
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 10186
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 10187
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 10188
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 10189
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 10190
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 10191
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 10192
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 10193
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 10194
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 10195
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 10196
,( 8, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 10197
,( 8, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 10198
,( 8, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 10199
,( 8, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 10200
,( 8, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 10201
,( 8, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 10202
,( 8, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 10203
,( 8, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 10204
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 10205
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 10206
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 10207
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 10208
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 10209
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 10210
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 10211
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 10212
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 10213
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 10214
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 10215
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 10216
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 10217
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 10218
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 10219
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 10220
,( 8, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 10221
,( 8, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 10222
,( 8, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 10223
,( 8, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 10224
,( 8, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 10225
,( 8, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 10226
,( 8, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 10227
,( 8, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 10228
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 10229
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 10230
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 10231
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 10232
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 10233
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 10234
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 10235
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 10236
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 10237
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 10238
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 10239
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 10240
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 10241
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 10242
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 10243
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 10244
,( 8, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 10245
,( 8, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 10246
,( 8, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 10247
,( 8, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 10248
,( 8, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 10249
,( 8, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 10250
,( 8, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 10251
,( 8, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 10252
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 10253
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 10254
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 10255
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 10256
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 10257
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 10258
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 10259
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 10260
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 10261
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 10262
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 10263
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 10264
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 10265
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 10266
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 10267
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 10268
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 10269
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 10270
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 10271
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 10272
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 10273
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 10274
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 10275
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 10276
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 16) -- 10277
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 16) -- 10278
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 16) -- 10279
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 16) -- 10280
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 16) -- 10281
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 16) -- 10282
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 16) -- 10283
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 16) -- 10284
,( 8, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 16) -- 10285
,( 8, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 16) -- 10286
,( 8, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 16) -- 10287
,( 8, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 16) -- 10288
,( 8, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 16) -- 10289
,( 8, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 16) -- 10290
,( 8, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 16) -- 10291
,( 8, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 16) -- 10292
,( 8, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 10293
,( 8, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 10294
,( 8, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 10295
,( 8, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 10296
,( 8, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 10297
,( 8, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 10298
,( 8, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 10299
,( 8, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 10300
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 16) -- 10301
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 16) -- 10302
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 16) -- 10303
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 16) -- 10304
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 16) -- 10305
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 16) -- 10306
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 16) -- 10307
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 16) -- 10308
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 16) -- 10309
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 16) -- 10310
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 16) -- 10311
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 16) -- 10312
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 16) -- 10313
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 16) -- 10314
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 16) -- 10315
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 16) -- 10316
,( 8, E,0,0,((28,28),(21,21),( 0, 0),(16,16),(18,18),(11,11)), 0, 15) -- 10317
,( 8, E,0,0,((29,29),(22,22),( 1, 1),(17,17),(19,19),(12,12)), 0, 15) -- 10318
,( 8, E,0,0,((30,30),(23,23),( 2, 2),(18,18),(20,20),(13,13)), 0, 15) -- 10319
,( 8, E,0,0,((31,31),(24,24),( 3, 3),(19,19),(21,21),(14,14)), 0, 15) -- 10320
,( 8, E,0,0,((32,32),(25,25),( 4, 4),(20,20),(22,22),(15,15)), 0, 15) -- 10321
,( 8, E,0,0,((33,33),(26,26),( 5, 5),(21,21),(23,23),(16,16)), 0, 15) -- 10322
,( 8, E,0,0,((34,34),(27,27),( 6, 6),(22,22),(24,24),(17,17)), 0, 15) -- 10323
,( 8, E,0,0,((35,35),(28,28),( 7, 7),(23,23),(25,25),(18,18)), 0, 15) -- 10324
,( 8, E,0,0,((28,28),(21,21),( 0, 0),(16,16),(18,18),(10,10)), 0, 15) -- 10325
,( 8, E,0,0,((29,29),(22,22),( 1, 1),(17,17),(19,19),(11,11)), 0, 15) -- 10326
,( 8, E,0,0,((30,30),(23,23),( 2, 2),(18,18),(20,20),(12,12)), 0, 15) -- 10327
,( 8, E,0,0,((31,31),(24,24),( 3, 3),(19,19),(21,21),(13,13)), 0, 15) -- 10328
,( 8, E,0,0,((32,32),(25,25),( 4, 4),(20,20),(22,22),(14,14)), 0, 15) -- 10329
,( 8, E,0,0,((33,33),(26,26),( 5, 5),(21,21),(23,23),(15,15)), 0, 15) -- 10330
,( 8, E,0,0,((34,34),(27,27),( 6, 6),(22,22),(24,24),(16,16)), 0, 15) -- 10331
,( 8, E,0,0,((35,35),(28,28),( 7, 7),(23,23),(25,25),(17,17)), 0, 15) -- 10332
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 10333
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 10334
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 10335
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 10336
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 10337
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 10338
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 10339
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 10340
,( 8, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 10341
,( 8, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 10342
,( 8, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 10343
,( 8, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 10344
,( 8, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 10345
,( 8, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 10346
,( 8, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 10347
,( 8, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 10348
,( 8, E,0,0,((26,29),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 14) -- 10349
,( 8, E,0,0,((28,31),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 14) -- 10350
,( 8, E,0,0,((30,33),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 14) -- 10351
,( 8, E,0,0,((32,35),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 14) -- 10352
,( 8, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(18,19),(10,13)), 0, 14) -- 10353
,( 8, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(20,21),(12,15)), 0, 14) -- 10354
,( 8, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(22,23),(14,17)), 0, 14) -- 10355
,( 8, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(24,25),(16,19)), 0, 14) -- 10356
,( 8, E,0,0,((26,29),(22,23),( 0, 1),(18,18),(20,21),(12,15)), 0, 14) -- 10357
,( 8, E,0,0,((28,31),(24,25),( 2, 3),(20,20),(22,23),(14,17)), 0, 14) -- 10358
,( 8, E,0,0,((30,33),(26,27),( 4, 5),(22,22),(24,25),(16,19)), 0, 14) -- 10359
,( 8, E,0,0,((32,35),(28,29),( 6, 7),(24,24),(26,27),(18,21)), 0, 14) -- 10360
,( 8, E,0,0,((26,29),(22,23),( 1, 1),(18,18),(19,19),(10,13)), 0, 13) -- 10361
,( 8, E,0,0,((28,31),(24,25),( 3, 3),(20,20),(21,21),(12,15)), 0, 13) -- 10362
,( 8, E,0,0,((30,33),(26,27),( 5, 5),(22,22),(23,23),(14,17)), 0, 13) -- 10363
,( 8, E,0,0,((32,35),(28,29),( 7, 7),(24,24),(25,25),(16,19)), 0, 13) -- 10364
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(17,17),(20,20),(12,15)), 0, 13) -- 10365
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(19,19),(22,22),(14,17)), 0, 13) -- 10366
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(21,21),(24,24),(16,19)), 0, 13) -- 10367
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(23,23),(26,26),(18,21)), 0, 13) -- 10368
,( 8, E,0,0,((26,29),(22,22),( 0, 1),(17,17),(20,20),(10,13)), 0, 13) -- 10369
,( 8, E,0,0,((28,31),(24,24),( 2, 3),(19,19),(22,22),(12,15)), 0, 13) -- 10370
,( 8, E,0,0,((30,33),(26,26),( 4, 5),(21,21),(24,24),(14,17)), 0, 13) -- 10371
,( 8, E,0,0,((32,35),(28,28),( 6, 7),(23,23),(26,26),(16,19)), 0, 13) -- 10372
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 10373
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 10374
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 10375
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 10376
,( 8, E,0,0,((26,29),(22,22),( 1, 1),(19,19),(20,21),(12,15)), 0, 12) -- 10377
,( 8, E,0,0,((28,31),(24,24),( 3, 3),(21,21),(22,23),(14,17)), 0, 12) -- 10378
,( 8, E,0,0,((30,33),(26,26),( 5, 5),(23,23),(24,25),(16,19)), 0, 12) -- 10379
,( 8, E,0,0,((32,35),(28,28),( 7, 7),(25,25),(26,27),(18,21)), 0, 12) -- 10380
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(16,17),(18,19),(10,13)), 0, 12) -- 10381
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(18,19),(20,21),(12,15)), 0, 12) -- 10382
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(20,21),(22,23),(14,17)), 0, 12) -- 10383
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(22,23),(24,25),(16,19)), 0, 12) -- 10384
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 12) -- 10385
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 12) -- 10386
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 12) -- 10387
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 12) -- 10388
,( 8, E,0,0,((26,29),(22,23),( 1, 1),(18,18),(20,20),(10,11)), 0, 12) -- 10389
,( 8, E,0,0,((28,31),(24,25),( 3, 3),(20,20),(22,22),(12,13)), 0, 12) -- 10390
,( 8, E,0,0,((30,33),(26,27),( 5, 5),(22,22),(24,24),(14,15)), 0, 12) -- 10391
,( 8, E,0,0,((32,35),(28,29),( 7, 7),(24,24),(26,26),(16,17)), 0, 12) -- 10392
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 10393
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 10394
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 10395
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 10396
,( 8, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(10,13)), 0, 11) -- 10397
,( 8, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(12,15)), 0, 11) -- 10398
,( 8, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(14,17)), 0, 11) -- 10399
,( 8, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(16,19)), 0, 11) -- 10400
,( 8, E,0,0,((22,25),(19,19),( 0, 0),(18,18),(20,21),(12,15)), 0, 11) -- 10401
,( 8, E,0,0,((24,27),(21,21),( 2, 2),(20,20),(22,23),(14,17)), 0, 11) -- 10402
,( 8, E,0,0,((26,29),(23,23),( 4, 4),(22,22),(24,25),(16,19)), 0, 11) -- 10403
,( 8, E,0,0,((28,31),(25,25),( 6, 6),(24,24),(26,27),(18,21)), 0, 11) -- 10404
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(16,17),(18,19),( 6, 9)), 0, 11) -- 10405
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(18,19),(20,21),( 8,11)), 0, 11) -- 10406
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(20,21),(22,23),(10,13)), 0, 11) -- 10407
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(22,23),(24,25),(12,15)), 0, 11) -- 10408
,( 8, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(20,21),(12,15)), 0, 11) -- 10409
,( 8, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(22,23),(14,17)), 0, 11) -- 10410
,( 8, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(24,25),(16,19)), 0, 11) -- 10411
,( 8, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(26,27),(18,21)), 0, 11) -- 10412
,( 8, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,22),(10,13)), 0, 10) -- 10413
,( 8, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,24),(12,15)), 0, 10) -- 10414
,( 8, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,26),(14,17)), 0, 10) -- 10415
,( 8, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,28),(16,19)), 0, 10) -- 10416
,( 8, E,0,0,((22,25),(18,19),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 10417
,( 8, E,0,0,((24,27),(20,21),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 10418
,( 8, E,0,0,((26,29),(22,23),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 10419
,( 8, E,0,0,((28,31),(24,25),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 10420
,( 8, E,0,0,((22,25),(18,19),( 0, 1),(18,19),(20,21),( 8,11)), 0, 10) -- 10421
,( 8, E,0,0,((24,27),(20,21),( 2, 3),(20,21),(22,23),(10,13)), 0, 10) -- 10422
,( 8, E,0,0,((26,29),(22,23),( 4, 5),(22,23),(24,25),(12,15)), 0, 10) -- 10423
,( 8, E,0,0,((28,31),(24,25),( 6, 7),(24,25),(26,27),(14,17)), 0, 10) -- 10424
,( 8, E,0,0,((22,25),(18,19),( 0, 0),(17,17),(20,20),( 8,11)), 0, 10) -- 10425
,( 8, E,0,0,((24,27),(20,21),( 2, 2),(19,19),(22,22),(10,13)), 0, 10) -- 10426
,( 8, E,0,0,((26,29),(22,23),( 4, 4),(21,21),(24,24),(12,15)), 0, 10) -- 10427
,( 8, E,0,0,((28,31),(24,25),( 6, 6),(23,23),(26,26),(14,17)), 0, 10) -- 10428
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(14,17)), 0, 10) -- 10429
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(16,19)), 0, 10) -- 10430
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(18,21)), 0, 10) -- 10431
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(20,23)), 0, 10) -- 10432
,( 8, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(12,15)), 0, 10) -- 10433
,( 8, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(14,17)), 0, 10) -- 10434
,( 8, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(16,19)), 0, 10) -- 10435
,( 8, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(18,21)), 0, 10) -- 10436
,( 8, E,0,0,((23,23),(20,20),( 1, 1),(18,19),(22,23),(12,15)), 0, 10) -- 10437
,( 8, E,0,0,((25,25),(22,22),( 3, 3),(20,21),(24,25),(14,17)), 0, 10) -- 10438
,( 8, E,0,0,((27,27),(24,24),( 5, 5),(22,23),(26,27),(16,19)), 0, 10) -- 10439
,( 8, E,0,0,((29,29),(26,26),( 7, 7),(24,25),(28,29),(18,21)), 0, 10) -- 10440
,( 8, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(21,21),(12,15)), 0, 10) -- 10441
,( 8, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(23,23),(14,17)), 0, 10) -- 10442
,( 8, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(25,25),(16,19)), 0, 10) -- 10443
,( 8, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(27,27),(18,21)), 0, 10) -- 10444
,( 8, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(18,19),( 8,11)), 0, 10) -- 10445
,( 8, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(20,21),(10,13)), 0, 10) -- 10446
,( 8, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(22,23),(12,15)), 0, 10) -- 10447
,( 8, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(24,25),(14,17)), 0, 10) -- 10448
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(10,13)), 0,  9) -- 10449
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(12,15)), 0,  9) -- 10450
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(14,17)), 0,  9) -- 10451
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(16,19)), 0,  9) -- 10452
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 10453
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 10454
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 10455
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 10456
,( 8, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 10457
,( 8, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 10458
,( 8, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 10459
,( 8, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 10460
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(20,21),(24,25),(14,17)), 0,  9) -- 10461
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(22,23),(26,27),(16,19)), 0,  9) -- 10462
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(24,25),(28,29),(18,21)), 0,  9) -- 10463
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(26,27),(30,31),(20,23)), 0,  9) -- 10464
,( 8, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 10465
,( 8, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 10466
,( 8, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 10467
,( 8, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 10468
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(18,19),( 4, 7)), 0,  9) -- 10469
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(20,21),( 6, 9)), 0,  9) -- 10470
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(22,23),( 8,11)), 0,  9) -- 10471
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(24,25),(10,13)), 0,  9) -- 10472
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 6, 9)), 0,  9) -- 10473
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),( 8,11)), 0,  9) -- 10474
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(10,13)), 0,  9) -- 10475
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(12,15)), 0,  9) -- 10476
,( 8, E,0,0,((18,21),(16,17),( 0, 0),(18,19),(20,21),( 6, 9)), 0,  9) -- 10477
,( 8, E,0,0,((20,23),(18,19),( 2, 2),(20,21),(22,23),( 8,11)), 0,  9) -- 10478
,( 8, E,0,0,((22,25),(20,21),( 4, 4),(22,23),(24,25),(10,13)), 0,  9) -- 10479
,( 8, E,0,0,((24,27),(22,23),( 6, 6),(24,25),(26,27),(12,15)), 0,  9) -- 10480
,( 8, E,0,0,((18,21),(16,17),( 0, 0),(18,19),(22,23),(10,13)), 0,  9) -- 10481
,( 8, E,0,0,((20,23),(18,19),( 2, 2),(20,21),(24,25),(12,15)), 0,  9) -- 10482
,( 8, E,0,0,((22,25),(20,21),( 4, 4),(22,23),(26,27),(14,17)), 0,  9) -- 10483
,( 8, E,0,0,((24,27),(22,23),( 6, 6),(24,25),(28,29),(16,19)), 0,  9) -- 10484
,( 8, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),(10,11)), 0,  9) -- 10485
,( 8, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),(12,13)), 0,  9) -- 10486
,( 8, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),(14,15)), 0,  9) -- 10487
,( 8, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),(16,17)), 0,  9) -- 10488
,( 8, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 6, 9)), 0,  9) -- 10489
,( 8, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 8,11)), 0,  9) -- 10490
,( 8, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),(10,13)), 0,  9) -- 10491
,( 8, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),(12,15)), 0,  9) -- 10492
,( 8, E,0,0,((23,23),(20,20),( 0, 1),(18,19),(20,21),(10,13)), 0,  9) -- 10493
,( 8, E,0,0,((25,25),(22,22),( 2, 3),(20,21),(22,23),(12,15)), 0,  9) -- 10494
,( 8, E,0,0,((27,27),(24,24),( 4, 5),(22,23),(24,25),(14,17)), 0,  9) -- 10495
,( 8, E,0,0,((29,29),(26,26),( 6, 7),(24,25),(26,27),(16,19)), 0,  9) -- 10496
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 10497
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 10498
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 10499
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 10500
,( 8, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(24,25),(16,19)), 0,  9) -- 10501
,( 8, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(26,27),(18,21)), 0,  9) -- 10502
,( 8, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(28,29),(20,23)), 0,  9) -- 10503
,( 8, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(30,31),(22,23)), 0,  9) -- 10504
,( 8, E,0,0,((23,23),(20,20),( 1, 1),(19,19),(22,22),( 8,11)), 0,  9) -- 10505
,( 8, E,0,0,((25,25),(22,22),( 3, 3),(21,21),(24,24),(10,13)), 0,  9) -- 10506
,( 8, E,0,0,((27,27),(24,24),( 5, 5),(23,23),(26,26),(12,15)), 0,  9) -- 10507
,( 8, E,0,0,((29,29),(26,26),( 7, 7),(25,25),(28,28),(14,17)), 0,  9) -- 10508
,( 8, E,0,0,((20,23),(18,19),( 0, 0),(17,17),(18,19),( 6, 9)), 0,  9) -- 10509
,( 8, E,0,0,((22,25),(20,21),( 2, 2),(19,19),(20,21),( 8,11)), 0,  9) -- 10510
,( 8, E,0,0,((24,27),(22,23),( 4, 4),(21,21),(22,23),(10,13)), 0,  9) -- 10511
,( 8, E,0,0,((26,29),(24,25),( 6, 6),(23,23),(24,25),(12,15)), 0,  9) -- 10512
,( 8, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(24,25),(10,13)), 0,  9) -- 10513
,( 8, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(26,27),(12,15)), 0,  9) -- 10514
,( 8, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(28,29),(14,17)), 0,  9) -- 10515
,( 8, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(30,31),(16,19)), 0,  9) -- 10516
,( 8, E,0,0,((22,25),(20,20),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 10517
,( 8, E,0,0,((24,27),(22,22),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 10518
,( 8, E,0,0,((26,29),(24,24),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 10519
,( 8, E,0,0,((28,31),(26,26),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 10520
,( 8, E,0,0,((18,21),(16,17),( 0, 0),(19,19),(24,25),(12,15)), 0,  9) -- 10521
,( 8, E,0,0,((20,23),(18,19),( 2, 2),(21,21),(26,27),(14,17)), 0,  9) -- 10522
,( 8, E,0,0,((22,25),(20,21),( 4, 4),(23,23),(28,29),(16,19)), 0,  9) -- 10523
,( 8, E,0,0,((24,27),(22,23),( 6, 6),(25,25),(30,31),(18,21)), 0,  9) -- 10524
,( 8, E,0,0,((20,23),(19,19),( 1, 1),(20,20),(22,23),( 6, 9)), 0,  9) -- 10525
,( 8, E,0,0,((22,25),(21,21),( 3, 3),(22,22),(24,25),( 8,11)), 0,  9) -- 10526
,( 8, E,0,0,((24,27),(23,23),( 5, 5),(24,24),(26,27),(10,13)), 0,  9) -- 10527
,( 8, E,0,0,((26,29),(25,25),( 7, 7),(26,26),(28,29),(12,15)), 0,  9) -- 10528
,( 8, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 10529
,( 8, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 10530
,( 8, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 10531
,( 8, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 10532
,( 8, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(22,25),( 8,11)), 0,  8) -- 10533
,( 8, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(24,27),(10,13)), 0,  8) -- 10534
,( 8, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(26,29),(12,15)), 0,  8) -- 10535
,( 8, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(28,31),(14,17)), 0,  8) -- 10536
,( 8, E,0,0,((18,21),(16,19),( 0, 1),(18,21),(18,21),(10,10)), 0,  8) -- 10537
,( 8, E,0,0,((20,23),(18,21),( 2, 3),(20,23),(20,23),(12,12)), 0,  8) -- 10538
,( 8, E,0,0,((22,25),(20,23),( 4, 5),(22,25),(22,25),(14,14)), 0,  8) -- 10539
,( 8, E,0,0,((24,27),(22,25),( 6, 7),(24,27),(24,27),(16,16)), 0,  8) -- 10540
,( 8, E,0,0,((14,17),(14,17),( 0, 1),(20,23),(24,27),(14,17)), 0,  8) -- 10541
,( 8, E,0,0,((16,19),(16,19),( 2, 3),(22,25),(26,29),(16,19)), 0,  8) -- 10542
,( 8, E,0,0,((18,21),(18,21),( 4, 5),(24,27),(28,31),(18,21)), 0,  8) -- 10543
,( 8, E,0,0,((20,23),(20,23),( 6, 7),(26,29),(30,33),(20,23)), 0,  8) -- 10544
,( 8, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(16,19),( 2, 5)), 0,  8) -- 10545
,( 8, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(18,21),( 4, 7)), 0,  8) -- 10546
,( 8, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(20,23),( 6, 9)), 0,  8) -- 10547
,( 8, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(22,25),( 8,11)), 0,  8) -- 10548
,( 8, E,0,0,((14,17),(14,17),( 0, 1),(18,21),(18,21),(99,99)), 0,  7) -- 10549
,( 8, E,0,0,((16,19),(16,19),( 2, 3),(20,23),(20,23),(99,99)), 0,  7) -- 10550
,( 8, E,0,0,((18,21),(18,21),( 4, 5),(22,25),(22,25),(99,99)), 0,  7) -- 10551
,( 8, E,0,0,((20,23),(20,23),( 6, 7),(24,27),(24,27),(99,99)), 0,  7) -- 10552
,( 8, E,0,0,((12,15),(14,17),( 0, 1),(18,21),(22,25),(99,99)), 0,  7) -- 10553
,( 8, E,0,0,((14,17),(16,19),( 2, 3),(20,23),(24,27),(99,99)), 0,  7) -- 10554
,( 8, E,0,0,((16,19),(18,21),( 4, 5),(22,25),(26,29),(99,99)), 0,  7) -- 10555
,( 8, E,0,0,((18,21),(20,23),( 6, 7),(24,27),(28,31),(99,99)), 0,  7) -- 10556
,( 8, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 10557
,( 8, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 10558
,( 8, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 10559
,( 8, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 10560
,( 8, E,0,1,((16,19),(16,19),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 10561
,( 8, E,0,1,((18,21),(18,21),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 10562
,( 8, E,0,1,((20,23),(20,23),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 10563
,( 8, E,0,1,((22,25),(22,25),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 10564
,( 8, E,0,1,((12,15),(12,15),( 0, 1),(20,23),(99,99),(99,99)), 0,  6) -- 10565
,( 8, E,0,1,((14,17),(14,17),( 2, 3),(22,25),(99,99),(99,99)), 0,  6) -- 10566
,( 8, E,0,1,((16,19),(16,19),( 4, 5),(24,27),(99,99),(99,99)), 0,  6) -- 10567
,( 8, E,0,1,((18,21),(18,21),( 6, 7),(26,29),(99,99),(99,99)), 0,  6) -- 10568
,( 8, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 10569
,( 8, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 10570
,( 8, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 10571
,( 8, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 10572
,( 8, E,0,1,((22,25),(20,23),( 0, 1),(13,13),(99,99),(99,99)), 0,  5) -- 10573
,( 8, E,0,1,((24,27),(22,25),( 2, 3),(15,15),(99,99),(99,99)), 0,  5) -- 10574
,( 8, E,0,1,((26,29),(24,27),( 4, 5),(17,17),(99,99),(99,99)), 0,  5) -- 10575
,( 8, E,0,1,((28,31),(26,29),( 6, 7),(19,19),(99,99),(99,99)), 0,  5) -- 10576
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 10577
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 10578
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 10579
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 10580
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 10581
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 10582
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 10583
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 10584
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 31) -- 10585
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 31) -- 10586
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 31) -- 10587
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(18,18),(10,10)), 1, 31) -- 10588
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(19,19),(11,11)), 1, 31) -- 10589
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(20,20),(12,12)), 1, 31) -- 10590
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(21,21),(13,13)), 1, 31) -- 10591
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(22,22),(14,14)), 1, 31) -- 10592
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 31) -- 10593
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 31) -- 10594
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 31) -- 10595
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 31) -- 10596
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 31) -- 10597
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 31) -- 10598
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 31) -- 10599
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 31) -- 10600
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 1, 31) -- 10601
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 1, 31) -- 10602
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 1, 31) -- 10603
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 1, 31) -- 10604
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 1, 31) -- 10605
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 1, 31) -- 10606
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 1, 31) -- 10607
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 1, 31) -- 10608
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 10609
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 10610
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 10611
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 10612
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 10613
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 10614
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 10615
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 10616
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 31) -- 10617
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 31) -- 10618
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 31) -- 10619
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 31) -- 10620
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 31) -- 10621
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 31) -- 10622
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 31) -- 10623
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 31) -- 10624
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 31) -- 10625
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 31) -- 10626
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(17,17),(10,10)), 1, 31) -- 10627
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(18,18),(11,11)), 1, 31) -- 10628
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(19,19),(12,12)), 1, 31) -- 10629
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(20,20),(13,13)), 1, 31) -- 10630
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(21,21),(14,14)), 1, 31) -- 10631
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(22,22),(15,15)), 1, 31) -- 10632
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 31) -- 10633
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 31) -- 10634
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 31) -- 10635
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 31) -- 10636
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 31) -- 10637
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 31) -- 10638
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 31) -- 10639
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 31) -- 10640
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 10641
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 10642
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 10643
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 10644
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 10645
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 10646
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 10647
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 10648
,( 9, E,0,0,((32,32),(23,23),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 30) -- 10649
,( 9, E,0,0,((33,33),(24,24),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 30) -- 10650
,( 9, E,0,0,((34,34),(25,25),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 30) -- 10651
,( 9, E,0,0,((35,35),(26,26),( 3, 3),(18,18),(18,18),(10,10)), 1, 30) -- 10652
,( 9, E,0,0,((36,36),(27,27),( 4, 4),(19,19),(19,19),(11,11)), 1, 30) -- 10653
,( 9, E,0,0,((37,37),(28,28),( 5, 5),(20,20),(20,20),(12,12)), 1, 30) -- 10654
,( 9, E,0,0,((38,38),(29,29),( 6, 6),(21,21),(21,21),(13,13)), 1, 30) -- 10655
,( 9, E,0,0,((39,39),(30,30),( 7, 7),(22,22),(22,22),(14,14)), 1, 30) -- 10656
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 28) -- 10657
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 28) -- 10658
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 28) -- 10659
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 28) -- 10660
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 28) -- 10661
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 28) -- 10662
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 28) -- 10663
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 28) -- 10664
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 27) -- 10665
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 27) -- 10666
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 27) -- 10667
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(18,18),(10,10)), 1, 27) -- 10668
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(19,19),(11,11)), 1, 27) -- 10669
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(20,20),(12,12)), 1, 27) -- 10670
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(21,21),(13,13)), 1, 27) -- 10671
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(22,22),(14,14)), 1, 27) -- 10672
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 26) -- 10673
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 26) -- 10674
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 26) -- 10675
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 26) -- 10676
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 26) -- 10677
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 26) -- 10678
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 26) -- 10679
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 26) -- 10680
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 25) -- 10681
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 25) -- 10682
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 25) -- 10683
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(18,18),(10,10)), 1, 25) -- 10684
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(19,19),(11,11)), 1, 25) -- 10685
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(20,20),(12,12)), 1, 25) -- 10686
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(21,21),(13,13)), 1, 25) -- 10687
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(22,22),(14,14)), 1, 25) -- 10688
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 25) -- 10689
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 25) -- 10690
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 25) -- 10691
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 25) -- 10692
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 25) -- 10693
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 25) -- 10694
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 25) -- 10695
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 25) -- 10696
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 24) -- 10697
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 24) -- 10698
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 24) -- 10699
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 24) -- 10700
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 24) -- 10701
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 24) -- 10702
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 24) -- 10703
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 24) -- 10704
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 10705
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 10706
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 10707
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 10708
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 10709
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 10710
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 10711
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 10712
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 24) -- 10713
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 24) -- 10714
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 24) -- 10715
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 24) -- 10716
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 24) -- 10717
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 24) -- 10718
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 24) -- 10719
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 24) -- 10720
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 23) -- 10721
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 23) -- 10722
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 23) -- 10723
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 23) -- 10724
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 23) -- 10725
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 23) -- 10726
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 23) -- 10727
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 23) -- 10728
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 22) -- 10729
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 22) -- 10730
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 22) -- 10731
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 22) -- 10732
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 22) -- 10733
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 22) -- 10734
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 22) -- 10735
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 22) -- 10736
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 21) -- 10737
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 21) -- 10738
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 21) -- 10739
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 21) -- 10740
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 21) -- 10741
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 21) -- 10742
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 21) -- 10743
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 21) -- 10744
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 21) -- 10745
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 21) -- 10746
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 21) -- 10747
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 21) -- 10748
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 21) -- 10749
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 21) -- 10750
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 21) -- 10751
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 21) -- 10752
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 21) -- 10753
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 21) -- 10754
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 21) -- 10755
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 21) -- 10756
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 21) -- 10757
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 21) -- 10758
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 21) -- 10759
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 21) -- 10760
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 20) -- 10761
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 20) -- 10762
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 20) -- 10763
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 20) -- 10764
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 20) -- 10765
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 20) -- 10766
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 20) -- 10767
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 20) -- 10768
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 20) -- 10769
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 20) -- 10770
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 20) -- 10771
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 20) -- 10772
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 20) -- 10773
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 20) -- 10774
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 20) -- 10775
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 20) -- 10776
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 10777
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 10778
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 10779
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 10780
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 10781
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 10782
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 10783
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 10784
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 10785
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 10786
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 10787
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 10788
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 10789
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 10790
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 10791
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 10792
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 19) -- 10793
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 19) -- 10794
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 19) -- 10795
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),(10,10)), 1, 19) -- 10796
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(11,11)), 1, 19) -- 10797
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(12,12)), 1, 19) -- 10798
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(13,13)), 1, 19) -- 10799
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(14,14)), 1, 19) -- 10800
,( 9, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 19) -- 10801
,( 9, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 19) -- 10802
,( 9, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 19) -- 10803
,( 9, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 19) -- 10804
,( 9, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 19) -- 10805
,( 9, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(10,10)), 1, 19) -- 10806
,( 9, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(11,11)), 1, 19) -- 10807
,( 9, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(12,12)), 1, 19) -- 10808
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 10809
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 10810
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 10811
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 10812
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 10813
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 10814
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 10815
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 10816
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 10817
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 10818
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 10819
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 10820
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 10821
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 10822
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 10823
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 10824
,( 9, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 10825
,( 9, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 10826
,( 9, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 10827
,( 9, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 10828
,( 9, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 10829
,( 9, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 10830
,( 9, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 10831
,( 9, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 10832
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 10833
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 10834
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 10835
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 10836
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 10837
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 10838
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 10839
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 10840
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 17) -- 10841
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 17) -- 10842
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 17) -- 10843
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 17) -- 10844
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 17) -- 10845
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 17) -- 10846
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 17) -- 10847
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 17) -- 10848
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 10849
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 10850
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 10851
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 10852
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 10853
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 10854
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 10855
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 10856
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 10857
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 10858
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 10859
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 10860
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 10861
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 10862
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 10863
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 10864
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 10865
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 10866
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 10867
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 10868
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 10869
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 10870
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 10871
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 10872
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 17) -- 10873
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 17) -- 10874
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 17) -- 10875
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 17) -- 10876
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 17) -- 10877
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 17) -- 10878
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 17) -- 10879
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 17) -- 10880
,( 9, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 10881
,( 9, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 10882
,( 9, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 10883
,( 9, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 10884
,( 9, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 10885
,( 9, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 10886
,( 9, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 10887
,( 9, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 10888
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 17) -- 10889
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 17) -- 10890
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 17) -- 10891
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 17) -- 10892
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 17) -- 10893
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 17) -- 10894
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 17) -- 10895
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 17) -- 10896
,( 9, E,0,0,((34,34),(24,24),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 10897
,( 9, E,0,0,((35,35),(25,25),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 10898
,( 9, E,0,0,((36,36),(26,26),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 10899
,( 9, E,0,0,((37,37),(27,27),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 10900
,( 9, E,0,0,((38,38),(28,28),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 10901
,( 9, E,0,0,((39,39),(29,29),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 10902
,( 9, E,0,0,((40,40),(30,30),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 10903
,( 9, E,0,0,((41,41),(31,31),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 10904
,( 9, E,0,0,((34,34),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 10905
,( 9, E,0,0,((35,35),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 10906
,( 9, E,0,0,((36,36),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 10907
,( 9, E,0,0,((37,37),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 10908
,( 9, E,0,0,((38,38),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 10909
,( 9, E,0,0,((39,39),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 10910
,( 9, E,0,0,((40,40),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 10911
,( 9, E,0,0,((41,41),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 10912
,( 9, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 10913
,( 9, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 10914
,( 9, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 10915
,( 9, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 10916
,( 9, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 10917
,( 9, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 10918
,( 9, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 10919
,( 9, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 10920
,( 9, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 16) -- 10921
,( 9, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 16) -- 10922
,( 9, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 16) -- 10923
,( 9, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 16) -- 10924
,( 9, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 16) -- 10925
,( 9, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 16) -- 10926
,( 9, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 16) -- 10927
,( 9, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 16) -- 10928
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 10929
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 10930
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 10931
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 10932
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 10933
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 10934
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 10935
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 10936
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 10937
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 10938
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 10939
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 10940
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 10941
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 10942
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 10943
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 10944
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 15) -- 10945
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 15) -- 10946
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 15) -- 10947
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 15) -- 10948
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 15) -- 10949
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(18,18),(10,10)), 1, 15) -- 10950
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(19,19),(11,11)), 1, 15) -- 10951
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(20,20),(12,12)), 1, 15) -- 10952
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 7, 7)), 1, 15) -- 10953
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 8, 8)), 1, 15) -- 10954
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 9, 9)), 1, 15) -- 10955
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),(10,10)), 1, 15) -- 10956
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(11,11)), 1, 15) -- 10957
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(12,12)), 1, 15) -- 10958
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(13,13)), 1, 15) -- 10959
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(14,14)), 1, 15) -- 10960
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(13,13),( 4, 4)), 1, 15) -- 10961
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(14,14),( 5, 5)), 1, 15) -- 10962
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(15,15),( 6, 6)), 1, 15) -- 10963
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(16,16),( 7, 7)), 1, 15) -- 10964
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(17,17),( 8, 8)), 1, 15) -- 10965
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(18,18),( 9, 9)), 1, 15) -- 10966
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(19,19),(10,10)), 1, 15) -- 10967
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(20,20),(11,11)), 1, 15) -- 10968
,( 9, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(13,13),( 4, 4)), 1, 15) -- 10969
,( 9, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(14,14),( 5, 5)), 1, 15) -- 10970
,( 9, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(15,15),( 6, 6)), 1, 15) -- 10971
,( 9, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(16,16),( 7, 7)), 1, 15) -- 10972
,( 9, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(17,17),( 8, 8)), 1, 15) -- 10973
,( 9, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(18,18),( 9, 9)), 1, 15) -- 10974
,( 9, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(19,19),(10,10)), 1, 15) -- 10975
,( 9, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(20,20),(11,11)), 1, 15) -- 10976
,( 9, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 15) -- 10977
,( 9, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 15) -- 10978
,( 9, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 15) -- 10979
,( 9, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 15) -- 10980
,( 9, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 15) -- 10981
,( 9, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 15) -- 10982
,( 9, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 15) -- 10983
,( 9, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 15) -- 10984
,( 9, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 10985
,( 9, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 10986
,( 9, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 10987
,( 9, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 10988
,( 9, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 10989
,( 9, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 10990
,( 9, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 10991
,( 9, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 10992
,( 9, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 10993
,( 9, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 10994
,( 9, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 10995
,( 9, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 10996
,( 9, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 10997
,( 9, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 10998
,( 9, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 10999
,( 9, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 11000
,( 9, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(13,13),( 5, 5)), 1, 15) -- 11001
,( 9, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(14,14),( 6, 6)), 1, 15) -- 11002
,( 9, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(15,15),( 7, 7)), 1, 15) -- 11003
,( 9, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(16,16),( 8, 8)), 1, 15) -- 11004
,( 9, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(17,17),( 9, 9)), 1, 15) -- 11005
,( 9, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(18,18),(10,10)), 1, 15) -- 11006
,( 9, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(19,19),(11,11)), 1, 15) -- 11007
,( 9, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(20,20),(12,12)), 1, 15) -- 11008
,( 9, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 11009
,( 9, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 11010
,( 9, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 11011
,( 9, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 11012
,( 9, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 11013
,( 9, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 11014
,( 9, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 11015
,( 9, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 11016
,( 9, E,0,0,((36,39),(26,27),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 11017
,( 9, E,0,0,((38,41),(28,29),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 11018
,( 9, E,0,0,((40,43),(30,31),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 11019
,( 9, E,0,0,((42,45),(32,33),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 11020
,( 9, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(13,13),( 4, 7)), 1, 13) -- 11021
,( 9, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(15,15),( 6, 9)), 1, 13) -- 11022
,( 9, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(17,17),( 8,11)), 1, 13) -- 11023
,( 9, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(19,19),(10,13)), 1, 13) -- 11024
,( 9, E,0,0,((38,38),(27,27),( 1, 1),(15,15),(14,14),( 4, 7)), 1, 13) -- 11025
,( 9, E,0,0,((40,40),(29,29),( 3, 3),(17,17),(16,16),( 6, 9)), 1, 13) -- 11026
,( 9, E,0,0,((42,42),(31,31),( 5, 5),(19,19),(18,18),( 8,11)), 1, 13) -- 11027
,( 9, E,0,0,((44,44),(33,33),( 7, 7),(21,21),(20,20),(10,13)), 1, 13) -- 11028
,( 9, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 11029
,( 9, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 11030
,( 9, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 11031
,( 9, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 11032
,( 9, E,0,0,((38,39),(27,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 11033
,( 9, E,0,0,((40,41),(29,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 11034
,( 9, E,0,0,((42,43),(31,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 11035
,( 9, E,0,0,((44,45),(33,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 11036
,( 9, E,0,0,((38,41),(28,29),( 1, 1),(15,15),(14,14),( 4, 7)), 1, 12) -- 11037
,( 9, E,0,0,((40,43),(30,31),( 3, 3),(17,17),(16,16),( 6, 9)), 1, 12) -- 11038
,( 9, E,0,0,((42,45),(32,33),( 5, 5),(19,19),(18,18),( 8,11)), 1, 12) -- 11039
,( 9, E,0,0,((44,47),(34,35),( 7, 7),(21,21),(20,20),(10,13)), 1, 12) -- 11040
,( 9, E,0,0,((38,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 12) -- 11041
,( 9, E,0,0,((40,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 12) -- 11042
,( 9, E,0,0,((42,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 12) -- 11043
,( 9, E,0,0,((44,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 12) -- 11044
,( 9, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 12) -- 11045
,( 9, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 12) -- 11046
,( 9, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 12) -- 11047
,( 9, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 12) -- 11048
,( 9, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 11049
,( 9, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 11050
,( 9, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 11051
,( 9, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 11052
,( 9, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(10,11),( 0, 3)), 1, 11) -- 11053
,( 9, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(12,13),( 2, 5)), 1, 11) -- 11054
,( 9, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(14,15),( 4, 7)), 1, 11) -- 11055
,( 9, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(16,17),( 6, 9)), 1, 11) -- 11056
,( 9, E,0,0,((38,41),(28,29),( 0, 1),(12,13),(10,11),( 0, 3)), 1, 11) -- 11057
,( 9, E,0,0,((40,43),(30,31),( 2, 3),(14,15),(12,13),( 2, 5)), 1, 11) -- 11058
,( 9, E,0,0,((42,45),(32,33),( 4, 5),(16,17),(14,15),( 4, 7)), 1, 11) -- 11059
,( 9, E,0,0,((44,47),(34,35),( 6, 7),(18,19),(16,17),( 6, 9)), 1, 11) -- 11060
,( 9, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 11) -- 11061
,( 9, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 11) -- 11062
,( 9, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 11) -- 11063
,( 9, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(18,18),( 8,11)), 1, 11) -- 11064
,( 9, E,0,0,((38,39),(27,27),( 0, 0),(14,14),(10,11),( 0, 3)), 1, 11) -- 11065
,( 9, E,0,0,((40,41),(29,29),( 2, 2),(16,16),(12,13),( 2, 5)), 1, 11) -- 11066
,( 9, E,0,0,((42,43),(31,31),( 4, 4),(18,18),(14,15),( 4, 7)), 1, 11) -- 11067
,( 9, E,0,0,((44,45),(33,33),( 6, 6),(20,20),(16,17),( 6, 9)), 1, 11) -- 11068
,( 9, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(10,11),( 4, 7)), 1, 10) -- 11069
,( 9, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(12,13),( 6, 9)), 1, 10) -- 11070
,( 9, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(14,15),( 8,11)), 1, 10) -- 11071
,( 9, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(16,17),(10,13)), 1, 10) -- 11072
,( 9, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 8,11)), 1, 10) -- 11073
,( 9, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(10,13)), 1, 10) -- 11074
,( 9, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(12,15)), 1, 10) -- 11075
,( 9, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(14,17)), 1, 10) -- 11076
,( 9, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 11077
,( 9, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 11078
,( 9, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 11079
,( 9, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 11080
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1, 10) -- 11081
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(10,11),( 2, 5)), 1, 10) -- 11082
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(12,13),( 4, 7)), 1, 10) -- 11083
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(14,15),( 6, 9)), 1, 10) -- 11084
,( 9, E,0,0,((42,42),(29,29),( 1, 1),(14,15),(12,13),( 4, 7)), 1, 10) -- 11085
,( 9, E,0,0,((44,44),(31,31),( 3, 3),(16,17),(14,15),( 6, 9)), 1, 10) -- 11086
,( 9, E,0,0,((46,46),(33,33),( 5, 5),(18,19),(16,17),( 8,11)), 1, 10) -- 11087
,( 9, E,0,0,((48,48),(35,35),( 7, 7),(20,21),(18,19),(10,13)), 1, 10) -- 11088
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(11,11),( 2, 5)), 1, 10) -- 11089
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(13,13),( 4, 7)), 1, 10) -- 11090
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(15,15),( 6, 9)), 1, 10) -- 11091
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(17,17),( 8,11)), 1, 10) -- 11092
,( 9, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(11,11),( 4, 5)), 1, 10) -- 11093
,( 9, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(13,13),( 6, 7)), 1, 10) -- 11094
,( 9, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(15,15),( 8, 9)), 1, 10) -- 11095
,( 9, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(17,17),(10,11)), 1, 10) -- 11096
,( 9, E,0,0,((38,41),(28,28),( 0, 0),(13,13),(12,12),( 4, 7)), 1, 10) -- 11097
,( 9, E,0,0,((40,43),(30,30),( 2, 2),(15,15),(14,14),( 6, 9)), 1, 10) -- 11098
,( 9, E,0,0,((42,45),(32,32),( 4, 4),(17,17),(16,16),( 8,11)), 1, 10) -- 11099
,( 9, E,0,0,((44,47),(34,34),( 6, 6),(19,19),(18,18),(10,13)), 1, 10) -- 11100
,( 9, E,0,0,((36,39),(26,27),( 0, 0),(14,14),(12,13),( 6, 9)), 1, 10) -- 11101
,( 9, E,0,0,((38,41),(28,29),( 2, 2),(16,16),(14,15),( 8,11)), 1, 10) -- 11102
,( 9, E,0,0,((40,43),(30,31),( 4, 4),(18,18),(16,17),(10,13)), 1, 10) -- 11103
,( 9, E,0,0,((42,45),(32,33),( 6, 6),(20,20),(18,19),(12,15)), 1, 10) -- 11104
,( 9, E,0,0,((42,45),(30,30),( 1, 1),(14,15),(12,13),( 4, 7)), 1, 10) -- 11105
,( 9, E,0,0,((44,47),(32,32),( 3, 3),(16,17),(14,15),( 6, 9)), 1, 10) -- 11106
,( 9, E,0,0,((46,49),(34,34),( 5, 5),(18,19),(16,17),( 8,11)), 1, 10) -- 11107
,( 9, E,0,0,((48,51),(36,36),( 7, 7),(20,21),(18,19),(10,13)), 1, 10) -- 11108
,( 9, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 11109
,( 9, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 11110
,( 9, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 11111
,( 9, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 11112
,( 9, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),( 8,11)), 1,  9) -- 11113
,( 9, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),(10,13)), 1,  9) -- 11114
,( 9, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(12,15)), 1,  9) -- 11115
,( 9, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(14,17)), 1,  9) -- 11116
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(13,13),(12,13),( 8,11)), 1,  9) -- 11117
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(15,15),(14,15),(10,13)), 1,  9) -- 11118
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(17,17),(16,17),(12,15)), 1,  9) -- 11119
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(19,19),(18,19),(14,17)), 1,  9) -- 11120
,( 9, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 2, 5)), 1,  9) -- 11121
,( 9, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 4, 7)), 1,  9) -- 11122
,( 9, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 6, 9)), 1,  9) -- 11123
,( 9, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 8,11)), 1,  9) -- 11124
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(12,13),( 8,11)), 1,  9) -- 11125
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(14,15),(10,13)), 1,  9) -- 11126
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(16,17),(12,15)), 1,  9) -- 11127
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(18,19),(14,17)), 1,  9) -- 11128
,( 9, E,0,0,((42,43),(29,29),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 11129
,( 9, E,0,0,((44,45),(31,31),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 11130
,( 9, E,0,0,((46,47),(33,33),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 11131
,( 9, E,0,0,((48,49),(35,35),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 11132
,( 9, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 11133
,( 9, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 11134
,( 9, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(10,13)), 1,  9) -- 11135
,( 9, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(12,15)), 1,  9) -- 11136
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(14,15),(12,15)), 1,  9) -- 11137
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(16,17),(14,17)), 1,  9) -- 11138
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(18,19),(16,19)), 1,  9) -- 11139
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(20,21),(18,21)), 1,  9) -- 11140
,( 9, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1,  9) -- 11141
,( 9, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 8,11)), 1,  9) -- 11142
,( 9, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(10,13)), 1,  9) -- 11143
,( 9, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(12,15)), 1,  9) -- 11144
,( 9, E,0,0,((42,45),(30,30),( 1, 1),(14,15),(14,15),(10,13)), 1,  9) -- 11145
,( 9, E,0,0,((44,47),(32,32),( 3, 3),(16,17),(16,17),(12,15)), 1,  9) -- 11146
,( 9, E,0,0,((46,49),(34,34),( 5, 5),(18,19),(18,19),(14,17)), 1,  9) -- 11147
,( 9, E,0,0,((48,51),(36,36),( 7, 7),(20,21),(20,21),(16,19)), 1,  9) -- 11148
,( 9, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,12),( 4, 7)), 1,  9) -- 11149
,( 9, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,14),( 6, 9)), 1,  9) -- 11150
,( 9, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,16),( 8,11)), 1,  9) -- 11151
,( 9, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,18),(10,13)), 1,  9) -- 11152
,( 9, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 6, 9)), 1,  9) -- 11153
,( 9, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 8,11)), 1,  9) -- 11154
,( 9, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),(10,13)), 1,  9) -- 11155
,( 9, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),(12,15)), 1,  9) -- 11156
,( 9, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),(10,10)), 1,  9) -- 11157
,( 9, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),(12,12)), 1,  9) -- 11158
,( 9, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(14,14)), 1,  9) -- 11159
,( 9, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(16,16)), 1,  9) -- 11160
,( 9, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),(12,15)), 1,  9) -- 11161
,( 9, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),(14,17)), 1,  9) -- 11162
,( 9, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(16,19)), 1,  9) -- 11163
,( 9, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(18,21)), 1,  9) -- 11164
,( 9, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 1)), 1,  9) -- 11165
,( 9, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 3)), 1,  9) -- 11166
,( 9, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 5)), 1,  9) -- 11167
,( 9, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 7)), 1,  9) -- 11168
,( 9, E,0,0,((42,45),(30,30),( 1, 1),(14,15),(13,13),(12,15)), 1,  9) -- 11169
,( 9, E,0,0,((44,47),(32,32),( 3, 3),(16,17),(15,15),(14,17)), 1,  9) -- 11170
,( 9, E,0,0,((46,49),(34,34),( 5, 5),(18,19),(17,17),(16,19)), 1,  9) -- 11171
,( 9, E,0,0,((48,51),(36,36),( 7, 7),(20,21),(19,19),(18,21)), 1,  9) -- 11172
,( 9, E,0,0,((46,49),(32,32),( 1, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 11173
,( 9, E,0,0,((48,51),(34,34),( 3, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 11174
,( 9, E,0,0,((50,53),(36,36),( 5, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 11175
,( 9, E,0,0,((52,55),(38,38),( 7, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 11176
,( 9, E,0,0,((40,43),(29,29),( 0, 0),(12,13),( 9, 9),( 4, 7)), 1,  9) -- 11177
,( 9, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(11,11),( 6, 9)), 1,  9) -- 11178
,( 9, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(13,13),( 8,11)), 1,  9) -- 11179
,( 9, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(15,15),(10,13)), 1,  9) -- 11180
,( 9, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(12,13),(12,15)), 1,  9) -- 11181
,( 9, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(14,15),(14,17)), 1,  9) -- 11182
,( 9, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(16,17),(16,19)), 1,  9) -- 11183
,( 9, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(18,19),(18,21)), 1,  9) -- 11184
,( 9, E,0,0,((44,47),(32,32),( 1, 1),(12,13),(11,11),( 9, 9)), 1,  9) -- 11185
,( 9, E,0,0,((46,49),(34,34),( 3, 3),(14,15),(13,13),(11,11)), 1,  9) -- 11186
,( 9, E,0,0,((48,51),(36,36),( 5, 5),(16,17),(15,15),(13,13)), 1,  9) -- 11187
,( 9, E,0,0,((50,53),(38,38),( 7, 7),(18,19),(17,17),(15,15)), 1,  9) -- 11188
,( 9, E,0,0,((42,42),(29,29),( 0, 0),(13,13),(10,10),( 0, 1)), 1,  9) -- 11189
,( 9, E,0,0,((44,44),(31,31),( 2, 2),(15,15),(12,12),( 2, 3)), 1,  9) -- 11190
,( 9, E,0,0,((46,46),(33,33),( 4, 4),(17,17),(14,14),( 4, 5)), 1,  9) -- 11191
,( 9, E,0,0,((48,48),(35,35),( 6, 6),(19,19),(16,16),( 6, 7)), 1,  9) -- 11192
,( 9, E,0,0,((42,42),(29,29),( 1, 1),(15,15),(14,14),( 8,11)), 1,  9) -- 11193
,( 9, E,0,0,((44,44),(31,31),( 3, 3),(17,17),(16,16),(10,13)), 1,  9) -- 11194
,( 9, E,0,0,((46,46),(33,33),( 5, 5),(19,19),(18,18),(12,15)), 1,  9) -- 11195
,( 9, E,0,0,((48,48),(35,35),( 7, 7),(21,21),(20,20),(14,17)), 1,  9) -- 11196
,( 9, E,0,0,((39,39),(27,27),( 0, 0),(13,13),(12,13),( 8,11)), 1,  9) -- 11197
,( 9, E,0,0,((41,41),(29,29),( 2, 2),(15,15),(14,15),(10,13)), 1,  9) -- 11198
,( 9, E,0,0,((43,43),(31,31),( 4, 4),(17,17),(16,17),(12,15)), 1,  9) -- 11199
,( 9, E,0,0,((45,45),(33,33),( 6, 6),(19,19),(18,19),(14,17)), 1,  9) -- 11200
,( 9, E,0,0,((44,47),(30,31),( 0, 1),(12,13),( 6, 7),(99,99)), 1,  9) -- 11201
,( 9, E,0,0,((46,49),(32,33),( 2, 3),(14,15),( 8, 9),(99,99)), 1,  9) -- 11202
,( 9, E,0,0,((48,51),(34,35),( 4, 5),(16,17),(10,11),(99,99)), 1,  9) -- 11203
,( 9, E,0,0,((50,53),(36,37),( 6, 7),(18,19),(12,13),(99,99)), 1,  9) -- 11204
,( 9, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(10,13),( 4, 7)), 1,  8) -- 11205
,( 9, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(12,15),( 6, 9)), 1,  8) -- 11206
,( 9, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(14,17),( 8,11)), 1,  8) -- 11207
,( 9, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(16,19),(10,13)), 1,  8) -- 11208
,( 9, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(16,16)), 1,  8) -- 11209
,( 9, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(18,18)), 1,  8) -- 11210
,( 9, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(20,20)), 1,  8) -- 11211
,( 9, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(22,22)), 1,  8) -- 11212
,( 9, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 8,11),(10,13)), 1,  8) -- 11213
,( 9, E,0,0,((46,49),(32,35),( 2, 3),(12,15),(10,13),(12,15)), 1,  8) -- 11214
,( 9, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(12,15),(14,17)), 1,  8) -- 11215
,( 9, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(14,17),(16,19)), 1,  8) -- 11216
,( 9, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(10,13),(10,13)), 1,  8) -- 11217
,( 9, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(12,15),(12,15)), 1,  8) -- 11218
,( 9, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(14,17),(14,17)), 1,  8) -- 11219
,( 9, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(16,19),(16,19)), 1,  8) -- 11220
,( 9, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  7) -- 11221
,( 9, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  7) -- 11222
,( 9, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  7) -- 11223
,( 9, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  7) -- 11224
,( 9, E,0,0,((48,51),(32,35),( 0, 1),(10,13),( 8,11),(99,99)), 1,  7) -- 11225
,( 9, E,0,0,((50,53),(34,37),( 2, 3),(12,15),(10,13),(99,99)), 1,  7) -- 11226
,( 9, E,0,0,((52,55),(36,39),( 4, 5),(14,17),(12,15),(99,99)), 1,  7) -- 11227
,( 9, E,0,0,((54,57),(38,41),( 6, 7),(16,19),(14,17),(99,99)), 1,  7) -- 11228
,( 9, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(18,21),(99,99)), 1,  7) -- 11229
,( 9, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(20,23),(99,99)), 1,  7) -- 11230
,( 9, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(22,25),(99,99)), 1,  7) -- 11231
,( 9, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(24,27),(99,99)), 1,  7) -- 11232
,( 9, E,0,1,((48,51),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 11233
,( 9, E,0,1,((50,53),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 11234
,( 9, E,0,1,((52,55),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 11235
,( 9, E,0,1,((54,57),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 11236
,( 9, E,0,1,((50,53),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  6) -- 11237
,( 9, E,0,1,((52,55),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  6) -- 11238
,( 9, E,0,1,((54,57),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  6) -- 11239
,( 9, E,0,1,((56,59),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  6) -- 11240
,( 9, E,0,1,((46,49),(30,33),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 11241
,( 9, E,0,1,((48,51),(32,35),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 11242
,( 9, E,0,1,((50,53),(34,37),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 11243
,( 9, E,0,1,((52,55),(36,39),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 11244
,( 9, E,0,1,((42,45),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 11245
,( 9, E,0,1,((44,47),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 11246
,( 9, E,0,1,((46,49),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 11247
,( 9, E,0,1,((48,51),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 11248
,( 9, E,0,1,((54,57),(34,37),( 0, 1),( 8,11),(99,99),(99,99)), 1,  6) -- 11249
,( 9, E,0,1,((56,59),(36,39),( 2, 3),(10,13),(99,99),(99,99)), 1,  6) -- 11250
,( 9, E,0,1,((58,61),(38,41),( 4, 5),(12,15),(99,99),(99,99)), 1,  6) -- 11251
,( 9, E,0,1,((60,63),(40,43),( 6, 7),(14,17),(99,99),(99,99)), 1,  6) -- 11252
,( 9, E,0,1,((46,49),(28,31),( 0, 1),(18,21),(99,99),(99,99)), 1,  5) -- 11253
,( 9, E,0,1,((48,51),(30,33),( 2, 3),(20,23),(99,99),(99,99)), 1,  5) -- 11254
,( 9, E,0,1,((50,53),(32,35),( 4, 5),(22,25),(99,99),(99,99)), 1,  5) -- 11255
,( 9, E,0,1,((52,55),(34,37),( 6, 7),(24,27),(99,99),(99,99)), 1,  5) -- 11256
,( 9, E,0,1,((38,41),(24,27),( 0, 1),(22,25),(99,99),(99,99)), 1,  5) -- 11257
,( 9, E,0,1,((40,43),(26,29),( 2, 3),(24,27),(99,99),(99,99)), 1,  5) -- 11258
,( 9, E,0,1,((42,45),(28,31),( 4, 5),(26,29),(99,99),(99,99)), 1,  5) -- 11259
,( 9, E,0,1,((44,47),(30,33),( 6, 7),(28,31),(99,99),(99,99)), 1,  5) -- 11260
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 11261
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 11262
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 11263
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 11264
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 11265
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 11266
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 11267
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 11268
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 11269
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 11270
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 11271
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 11272
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 11273
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 11274
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 11275
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 11276
,( 9, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 11277
,( 9, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 11278
,( 9, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 11279
,( 9, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 11280
,( 9, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 11281
,( 9, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 11282
,( 9, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 11283
,( 9, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 11284
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 11285
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 11286
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 11287
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 11288
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 11289
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 11290
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 11291
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 11292
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 11293
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 11294
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 11295
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 11296
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 11297
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 11298
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 11299
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 11300
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 11301
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 11302
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 11303
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 11304
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 11305
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 11306
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 11307
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 11308
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(15,15),( 8, 8)), 0, 31) -- 11309
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(16,16),( 9, 9)), 0, 31) -- 11310
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(17,17),(10,10)), 0, 31) -- 11311
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(18,18),(11,11)), 0, 31) -- 11312
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(19,19),(12,12)), 0, 31) -- 11313
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(20,20),(13,13)), 0, 31) -- 11314
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(21,21),(14,14)), 0, 31) -- 11315
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(22,22),(15,15)), 0, 31) -- 11316
,( 9, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 30) -- 11317
,( 9, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 30) -- 11318
,( 9, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 30) -- 11319
,( 9, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 30) -- 11320
,( 9, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 30) -- 11321
,( 9, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 30) -- 11322
,( 9, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 30) -- 11323
,( 9, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 30) -- 11324
,( 9, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 29) -- 11325
,( 9, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 29) -- 11326
,( 9, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 29) -- 11327
,( 9, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 29) -- 11328
,( 9, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 29) -- 11329
,( 9, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 29) -- 11330
,( 9, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 29) -- 11331
,( 9, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 29) -- 11332
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 28) -- 11333
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 28) -- 11334
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 28) -- 11335
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 28) -- 11336
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 28) -- 11337
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 28) -- 11338
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 28) -- 11339
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 28) -- 11340
,( 9, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 27) -- 11341
,( 9, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 27) -- 11342
,( 9, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 27) -- 11343
,( 9, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 27) -- 11344
,( 9, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 27) -- 11345
,( 9, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 27) -- 11346
,( 9, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 27) -- 11347
,( 9, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 27) -- 11348
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 25) -- 11349
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 25) -- 11350
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 25) -- 11351
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 25) -- 11352
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 25) -- 11353
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 25) -- 11354
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 25) -- 11355
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 25) -- 11356
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 25) -- 11357
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 25) -- 11358
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 25) -- 11359
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 25) -- 11360
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 25) -- 11361
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 25) -- 11362
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 25) -- 11363
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 25) -- 11364
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 24) -- 11365
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 24) -- 11366
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 24) -- 11367
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 24) -- 11368
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 24) -- 11369
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 24) -- 11370
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 24) -- 11371
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 24) -- 11372
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 23) -- 11373
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 23) -- 11374
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 23) -- 11375
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 23) -- 11376
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 23) -- 11377
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 23) -- 11378
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 23) -- 11379
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 23) -- 11380
,( 9, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 23) -- 11381
,( 9, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 23) -- 11382
,( 9, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 23) -- 11383
,( 9, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 23) -- 11384
,( 9, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 23) -- 11385
,( 9, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 23) -- 11386
,( 9, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 23) -- 11387
,( 9, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 23) -- 11388
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 22) -- 11389
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 22) -- 11390
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 22) -- 11391
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 22) -- 11392
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 22) -- 11393
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 22) -- 11394
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 22) -- 11395
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 22) -- 11396
,( 9, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 11397
,( 9, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 11398
,( 9, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 11399
,( 9, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 11400
,( 9, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 11401
,( 9, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 11402
,( 9, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 11403
,( 9, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 11404
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 20) -- 11405
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 20) -- 11406
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 20) -- 11407
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 20) -- 11408
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 20) -- 11409
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 20) -- 11410
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 20) -- 11411
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 20) -- 11412
,( 9, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 20) -- 11413
,( 9, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(17,17),(10,10)), 0, 20) -- 11414
,( 9, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(18,18),(11,11)), 0, 20) -- 11415
,( 9, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(19,19),(12,12)), 0, 20) -- 11416
,( 9, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(20,20),(13,13)), 0, 20) -- 11417
,( 9, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(21,21),(14,14)), 0, 20) -- 11418
,( 9, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(22,22),(15,15)), 0, 20) -- 11419
,( 9, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(23,23),(16,16)), 0, 20) -- 11420
,( 9, E,0,0,((30,30),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 11421
,( 9, E,0,0,((31,31),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 11422
,( 9, E,0,0,((32,32),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 11423
,( 9, E,0,0,((33,33),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 11424
,( 9, E,0,0,((34,34),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 11425
,( 9, E,0,0,((35,35),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 11426
,( 9, E,0,0,((36,36),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 11427
,( 9, E,0,0,((37,37),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 11428
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(17,17),(10,10)), 0, 19) -- 11429
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(18,18),(11,11)), 0, 19) -- 11430
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(19,19),(12,12)), 0, 19) -- 11431
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(20,20),(13,13)), 0, 19) -- 11432
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(21,21),(14,14)), 0, 19) -- 11433
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(22,22),(15,15)), 0, 19) -- 11434
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(23,23),(16,16)), 0, 19) -- 11435
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(24,24),(17,17)), 0, 19) -- 11436
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 11437
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 11438
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 11439
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 11440
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 11441
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 11442
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 11443
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 11444
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 11445
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 11446
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 11447
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 11448
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 11449
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 11450
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 11451
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 11452
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 11453
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 11454
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 11455
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 11456
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 11457
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 11458
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 11459
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 11460
,( 9, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 11461
,( 9, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 11462
,( 9, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 11463
,( 9, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 11464
,( 9, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 11465
,( 9, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 11466
,( 9, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 11467
,( 9, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 11468
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 11469
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 11470
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 11471
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 11472
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 11473
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 11474
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 11475
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 11476
,( 9, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 11477
,( 9, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 11478
,( 9, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 11479
,( 9, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 11480
,( 9, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 11481
,( 9, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 11482
,( 9, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 11483
,( 9, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 11484
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 11485
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 11486
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 11487
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 11488
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 11489
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 11490
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 11491
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 11492
,( 9, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 11493
,( 9, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 11494
,( 9, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 11495
,( 9, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 11496
,( 9, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 11497
,( 9, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 11498
,( 9, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 11499
,( 9, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 11500
,( 9, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 11501
,( 9, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 11502
,( 9, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 11503
,( 9, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 11504
,( 9, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 11505
,( 9, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 11506
,( 9, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 11507
,( 9, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 11508
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 11509
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 11510
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 11511
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 11512
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 11513
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 11514
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 11515
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 11516
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 11517
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 11518
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 11519
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 11520
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 11521
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 11522
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 11523
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 11524
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 17) -- 11525
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 17) -- 11526
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 17) -- 11527
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 17) -- 11528
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 17) -- 11529
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 17) -- 11530
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 17) -- 11531
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 17) -- 11532
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(11,11)), 0, 17) -- 11533
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(12,12)), 0, 17) -- 11534
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(13,13)), 0, 17) -- 11535
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(14,14)), 0, 17) -- 11536
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(15,15)), 0, 17) -- 11537
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(16,16)), 0, 17) -- 11538
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(17,17)), 0, 17) -- 11539
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(18,18)), 0, 17) -- 11540
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(10,10)), 0, 16) -- 11541
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(11,11)), 0, 16) -- 11542
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(12,12)), 0, 16) -- 11543
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(13,13)), 0, 16) -- 11544
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(14,14)), 0, 16) -- 11545
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(15,15)), 0, 16) -- 11546
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(16,16)), 0, 16) -- 11547
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(17,17)), 0, 16) -- 11548
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 11549
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 11550
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 11551
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 11552
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 11553
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 11554
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 11555
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 11556
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 11557
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 11558
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 11559
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 11560
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 11561
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 11562
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 11563
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 11564
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 16) -- 11565
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 16) -- 11566
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 16) -- 11567
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 16) -- 11568
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 16) -- 11569
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 16) -- 11570
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 16) -- 11571
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 16) -- 11572
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 11573
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 11574
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 11575
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 11576
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 11577
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 11578
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 11579
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 11580
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 11581
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 11582
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 11583
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 11584
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 11585
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 11586
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 11587
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 11588
,( 9, E,0,0,((28,28),(21,21),( 0, 0),(16,16),(18,18),(11,11)), 0, 15) -- 11589
,( 9, E,0,0,((29,29),(22,22),( 1, 1),(17,17),(19,19),(12,12)), 0, 15) -- 11590
,( 9, E,0,0,((30,30),(23,23),( 2, 2),(18,18),(20,20),(13,13)), 0, 15) -- 11591
,( 9, E,0,0,((31,31),(24,24),( 3, 3),(19,19),(21,21),(14,14)), 0, 15) -- 11592
,( 9, E,0,0,((32,32),(25,25),( 4, 4),(20,20),(22,22),(15,15)), 0, 15) -- 11593
,( 9, E,0,0,((33,33),(26,26),( 5, 5),(21,21),(23,23),(16,16)), 0, 15) -- 11594
,( 9, E,0,0,((34,34),(27,27),( 6, 6),(22,22),(24,24),(17,17)), 0, 15) -- 11595
,( 9, E,0,0,((35,35),(28,28),( 7, 7),(23,23),(25,25),(18,18)), 0, 15) -- 11596
,( 9, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 11597
,( 9, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 11598
,( 9, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 11599
,( 9, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 11600
,( 9, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 11601
,( 9, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 11602
,( 9, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 11603
,( 9, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 11604
,( 9, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(10,10)), 0, 15) -- 11605
,( 9, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(11,11)), 0, 15) -- 11606
,( 9, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(12,12)), 0, 15) -- 11607
,( 9, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(13,13)), 0, 15) -- 11608
,( 9, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(14,14)), 0, 15) -- 11609
,( 9, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(15,15)), 0, 15) -- 11610
,( 9, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(16,16)), 0, 15) -- 11611
,( 9, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(17,17)), 0, 15) -- 11612
,( 9, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 11613
,( 9, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 11614
,( 9, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 11615
,( 9, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 11616
,( 9, E,0,0,((26,29),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 14) -- 11617
,( 9, E,0,0,((28,31),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 14) -- 11618
,( 9, E,0,0,((30,33),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 14) -- 11619
,( 9, E,0,0,((32,35),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 14) -- 11620
,( 9, E,0,0,((28,31),(22,23),( 1, 1),(18,18),(20,20),(12,15)), 0, 14) -- 11621
,( 9, E,0,0,((30,33),(24,25),( 3, 3),(20,20),(22,22),(14,17)), 0, 14) -- 11622
,( 9, E,0,0,((32,35),(26,27),( 5, 5),(22,22),(24,24),(16,19)), 0, 14) -- 11623
,( 9, E,0,0,((34,37),(28,29),( 7, 7),(24,24),(26,26),(18,21)), 0, 14) -- 11624
,( 9, E,0,0,((26,29),(22,23),( 0, 1),(18,18),(19,19),(10,13)), 0, 13) -- 11625
,( 9, E,0,0,((28,31),(24,25),( 2, 3),(20,20),(21,21),(12,15)), 0, 13) -- 11626
,( 9, E,0,0,((30,33),(26,27),( 4, 5),(22,22),(23,23),(14,17)), 0, 13) -- 11627
,( 9, E,0,0,((32,35),(28,29),( 6, 7),(24,24),(25,25),(16,19)), 0, 13) -- 11628
,( 9, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(12,15)), 0, 13) -- 11629
,( 9, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(14,17)), 0, 13) -- 11630
,( 9, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(16,19)), 0, 13) -- 11631
,( 9, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(18,21)), 0, 13) -- 11632
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 11633
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 11634
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 11635
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 11636
,( 9, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(12,15)), 0, 12) -- 11637
,( 9, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(14,17)), 0, 12) -- 11638
,( 9, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(16,19)), 0, 12) -- 11639
,( 9, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(18,21)), 0, 12) -- 11640
,( 9, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(18,19),(10,13)), 0, 12) -- 11641
,( 9, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(20,21),(12,15)), 0, 12) -- 11642
,( 9, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(22,23),(14,17)), 0, 12) -- 11643
,( 9, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(24,25),(16,19)), 0, 12) -- 11644
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 11645
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 11646
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 11647
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 11648
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 11649
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 11650
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 11651
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 11652
,( 9, E,0,0,((22,25),(19,19),( 0, 0),(18,18),(20,21),(12,15)), 0, 11) -- 11653
,( 9, E,0,0,((24,27),(21,21),( 2, 2),(20,20),(22,23),(14,17)), 0, 11) -- 11654
,( 9, E,0,0,((26,29),(23,23),( 4, 4),(22,22),(24,25),(16,19)), 0, 11) -- 11655
,( 9, E,0,0,((28,31),(25,25),( 6, 6),(24,24),(26,27),(18,21)), 0, 11) -- 11656
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(16,17),(18,19),( 8,11)), 0, 11) -- 11657
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(18,19),(20,21),(10,13)), 0, 11) -- 11658
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(20,21),(22,23),(12,15)), 0, 11) -- 11659
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(22,23),(24,25),(14,17)), 0, 11) -- 11660
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(18,18),(19,19),(10,13)), 0, 11) -- 11661
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(20,20),(21,21),(12,15)), 0, 11) -- 11662
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(22,22),(23,23),(14,17)), 0, 11) -- 11663
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(24,24),(25,25),(16,19)), 0, 11) -- 11664
,( 9, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 11665
,( 9, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 11666
,( 9, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 11667
,( 9, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 11668
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(14,17)), 0, 10) -- 11669
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(16,19)), 0, 10) -- 11670
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(18,21)), 0, 10) -- 11671
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(20,23)), 0, 10) -- 11672
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 8,11)), 0, 10) -- 11673
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),(10,13)), 0, 10) -- 11674
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(12,15)), 0, 10) -- 11675
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(14,17)), 0, 10) -- 11676
,( 9, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(18,19),( 6, 9)), 0, 10) -- 11677
,( 9, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(20,21),( 8,11)), 0, 10) -- 11678
,( 9, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(22,23),(10,13)), 0, 10) -- 11679
,( 9, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(24,25),(12,15)), 0, 10) -- 11680
,( 9, E,0,0,((23,23),(20,20),( 0, 1),(18,19),(20,21),(10,13)), 0, 10) -- 11681
,( 9, E,0,0,((25,25),(22,22),( 2, 3),(20,21),(22,23),(12,15)), 0, 10) -- 11682
,( 9, E,0,0,((27,27),(24,24),( 4, 5),(22,23),(24,25),(14,17)), 0, 10) -- 11683
,( 9, E,0,0,((29,29),(26,26),( 6, 7),(24,25),(26,27),(16,19)), 0, 10) -- 11684
,( 9, E,0,0,((22,25),(18,19),( 0, 0),(17,17),(20,21),(10,13)), 0, 10) -- 11685
,( 9, E,0,0,((24,27),(20,21),( 2, 2),(19,19),(22,23),(12,15)), 0, 10) -- 11686
,( 9, E,0,0,((26,29),(22,23),( 4, 4),(21,21),(24,25),(14,17)), 0, 10) -- 11687
,( 9, E,0,0,((28,31),(24,25),( 6, 6),(23,23),(26,27),(16,19)), 0, 10) -- 11688
,( 9, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(14,17)), 0, 10) -- 11689
,( 9, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(16,19)), 0, 10) -- 11690
,( 9, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(18,21)), 0, 10) -- 11691
,( 9, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(20,23)), 0, 10) -- 11692
,( 9, E,0,0,((24,25),(20,20),( 0, 0),(17,17),(20,20),( 8,11)), 0, 10) -- 11693
,( 9, E,0,0,((26,27),(22,22),( 2, 2),(19,19),(22,22),(10,13)), 0, 10) -- 11694
,( 9, E,0,0,((28,29),(24,24),( 4, 4),(21,21),(24,24),(12,15)), 0, 10) -- 11695
,( 9, E,0,0,((30,31),(26,26),( 6, 6),(23,23),(26,26),(14,17)), 0, 10) -- 11696
,( 9, E,0,0,((26,27),(22,22),( 1, 1),(18,19),(20,21),( 8,11)), 0, 10) -- 11697
,( 9, E,0,0,((28,29),(24,24),( 3, 3),(20,21),(22,23),(10,13)), 0, 10) -- 11698
,( 9, E,0,0,((30,31),(26,26),( 5, 5),(22,23),(24,25),(12,15)), 0, 10) -- 11699
,( 9, E,0,0,((32,33),(28,28),( 7, 7),(24,25),(26,27),(14,17)), 0, 10) -- 11700
,( 9, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(19,19),( 6, 9)), 0, 10) -- 11701
,( 9, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(21,21),( 8,11)), 0, 10) -- 11702
,( 9, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(23,23),(10,13)), 0, 10) -- 11703
,( 9, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(25,25),(12,15)), 0, 10) -- 11704
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(10,13)), 0,  9) -- 11705
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(12,15)), 0,  9) -- 11706
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(14,17)), 0,  9) -- 11707
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(16,19)), 0,  9) -- 11708
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(18,19),( 4, 7)), 0,  9) -- 11709
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(20,21),( 6, 9)), 0,  9) -- 11710
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(22,23),( 8,11)), 0,  9) -- 11711
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(24,25),(10,13)), 0,  9) -- 11712
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(20,20),(22,23),(10,13)), 0,  9) -- 11713
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(22,22),(24,25),(12,15)), 0,  9) -- 11714
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(24,24),(26,27),(14,17)), 0,  9) -- 11715
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(26,26),(28,29),(16,19)), 0,  9) -- 11716
,( 9, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 11717
,( 9, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 11718
,( 9, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 11719
,( 9, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 11720
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 4, 7)), 0,  9) -- 11721
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 6, 9)), 0,  9) -- 11722
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),( 8,11)), 0,  9) -- 11723
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(10,13)), 0,  9) -- 11724
,( 9, E,0,0,((20,23),(18,19),( 1, 1),(20,21),(24,25),(14,17)), 0,  9) -- 11725
,( 9, E,0,0,((22,25),(20,21),( 3, 3),(22,23),(26,27),(16,19)), 0,  9) -- 11726
,( 9, E,0,0,((24,27),(22,23),( 5, 5),(24,25),(28,29),(18,21)), 0,  9) -- 11727
,( 9, E,0,0,((26,29),(24,25),( 7, 7),(26,27),(30,31),(20,23)), 0,  9) -- 11728
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(21,21),(12,15)), 0,  9) -- 11729
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(23,23),(14,17)), 0,  9) -- 11730
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(25,25),(16,19)), 0,  9) -- 11731
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(27,27),(18,21)), 0,  9) -- 11732
,( 9, E,0,0,((18,21),(17,17),( 0, 0),(18,19),(22,23),(10,13)), 0,  9) -- 11733
,( 9, E,0,0,((20,23),(19,19),( 2, 2),(20,21),(24,25),(12,15)), 0,  9) -- 11734
,( 9, E,0,0,((22,25),(21,21),( 4, 4),(22,23),(26,27),(14,17)), 0,  9) -- 11735
,( 9, E,0,0,((24,27),(23,23),( 6, 6),(24,25),(28,29),(16,19)), 0,  9) -- 11736
,( 9, E,0,0,((22,25),(20,21),( 1, 1),(19,19),(22,23),( 8,11)), 0,  9) -- 11737
,( 9, E,0,0,((24,27),(22,23),( 3, 3),(21,21),(24,25),(10,13)), 0,  9) -- 11738
,( 9, E,0,0,((26,29),(24,25),( 5, 5),(23,23),(26,27),(12,15)), 0,  9) -- 11739
,( 9, E,0,0,((28,31),(26,27),( 7, 7),(25,25),(28,29),(14,17)), 0,  9) -- 11740
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 6, 9)), 0,  9) -- 11741
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),( 8,11)), 0,  9) -- 11742
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(10,13)), 0,  9) -- 11743
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(12,15)), 0,  9) -- 11744
,( 9, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 11745
,( 9, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 11746
,( 9, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 11747
,( 9, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 11748
,( 9, E,0,0,((18,21),(17,17),( 0, 1),(18,19),(20,21),( 4, 7)), 0,  9) -- 11749
,( 9, E,0,0,((20,23),(19,19),( 2, 3),(20,21),(22,23),( 6, 9)), 0,  9) -- 11750
,( 9, E,0,0,((22,25),(21,21),( 4, 5),(22,23),(24,25),( 8,11)), 0,  9) -- 11751
,( 9, E,0,0,((24,27),(23,23),( 6, 7),(24,25),(26,27),(10,13)), 0,  9) -- 11752
,( 9, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 11753
,( 9, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 11754
,( 9, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 11755
,( 9, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 11756
,( 9, E,0,0,((16,19),(16,17),( 0, 1),(20,21),(24,25),(16,19)), 0,  9) -- 11757
,( 9, E,0,0,((18,21),(18,19),( 2, 3),(22,23),(26,27),(18,21)), 0,  9) -- 11758
,( 9, E,0,0,((20,23),(20,21),( 4, 5),(24,25),(28,29),(20,23)), 0,  9) -- 11759
,( 9, E,0,0,((22,25),(22,23),( 6, 7),(26,27),(30,31),(22,23)), 0,  9) -- 11760
,( 9, E,0,0,((20,23),(18,19),( 0, 0),(17,17),(18,19),( 4, 7)), 0,  9) -- 11761
,( 9, E,0,0,((22,25),(20,21),( 2, 2),(19,19),(20,21),( 6, 9)), 0,  9) -- 11762
,( 9, E,0,0,((24,27),(22,23),( 4, 4),(21,21),(22,23),( 8,11)), 0,  9) -- 11763
,( 9, E,0,0,((26,29),(24,25),( 6, 6),(23,23),(24,25),(10,13)), 0,  9) -- 11764
,( 9, E,0,0,((22,25),(20,20),( 1, 1),(20,20),(24,24),(14,17)), 0,  9) -- 11765
,( 9, E,0,0,((24,27),(22,22),( 3, 3),(22,22),(26,26),(16,19)), 0,  9) -- 11766
,( 9, E,0,0,((26,29),(24,24),( 5, 5),(24,24),(28,28),(18,21)), 0,  9) -- 11767
,( 9, E,0,0,((28,31),(26,26),( 7, 7),(26,26),(30,30),(20,23)), 0,  9) -- 11768
,( 9, E,0,0,((22,25),(20,21),( 1, 1),(19,19),(20,21),( 2, 5)), 0,  9) -- 11769
,( 9, E,0,0,((24,27),(22,23),( 3, 3),(21,21),(22,23),( 4, 7)), 0,  9) -- 11770
,( 9, E,0,0,((26,29),(24,25),( 5, 5),(23,23),(24,25),( 6, 9)), 0,  9) -- 11771
,( 9, E,0,0,((28,31),(26,27),( 7, 7),(25,25),(26,27),( 8,11)), 0,  9) -- 11772
,( 9, E,0,0,((20,21),(18,19),( 1, 1),(20,21),(26,26),(16,19)), 0,  9) -- 11773
,( 9, E,0,0,((22,23),(20,21),( 3, 3),(22,23),(28,28),(18,21)), 0,  9) -- 11774
,( 9, E,0,0,((24,25),(22,23),( 5, 5),(24,25),(30,30),(20,23)), 0,  9) -- 11775
,( 9, E,0,0,((26,27),(24,25),( 7, 7),(26,27),(32,32),(22,23)), 0,  9) -- 11776
,( 9, E,0,0,((16,19),(16,17),( 0, 0),(18,19),(22,23),( 6, 9)), 0,  9) -- 11777
,( 9, E,0,0,((18,21),(18,19),( 2, 2),(20,21),(24,25),( 8,11)), 0,  9) -- 11778
,( 9, E,0,0,((20,23),(20,21),( 4, 4),(22,23),(26,27),(10,13)), 0,  9) -- 11779
,( 9, E,0,0,((22,25),(22,23),( 6, 6),(24,25),(28,29),(12,15)), 0,  9) -- 11780
,( 9, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(24,25),(10,13)), 0,  9) -- 11781
,( 9, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(26,27),(12,15)), 0,  9) -- 11782
,( 9, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(28,29),(14,17)), 0,  9) -- 11783
,( 9, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(30,31),(16,19)), 0,  9) -- 11784
,( 9, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(23,23),(14,14)), 0,  9) -- 11785
,( 9, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(25,25),(16,16)), 0,  9) -- 11786
,( 9, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(27,27),(18,18)), 0,  9) -- 11787
,( 9, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(29,29),(20,20)), 0,  9) -- 11788
,( 9, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 0, 3)), 0,  9) -- 11789
,( 9, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 2, 5)), 0,  9) -- 11790
,( 9, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),( 4, 7)), 0,  9) -- 11791
,( 9, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),( 6, 9)), 0,  9) -- 11792
,( 9, E,0,0,((18,21),(18,18),( 1, 1),(20,20),(22,23),( 6, 9)), 0,  9) -- 11793
,( 9, E,0,0,((20,23),(20,20),( 3, 3),(22,22),(24,25),( 8,11)), 0,  9) -- 11794
,( 9, E,0,0,((22,25),(22,22),( 5, 5),(24,24),(26,27),(10,13)), 0,  9) -- 11795
,( 9, E,0,0,((24,27),(24,24),( 7, 7),(26,26),(28,29),(12,15)), 0,  9) -- 11796
,( 9, E,0,0,((18,21),(16,19),( 0, 1),(18,21),(18,21),(10,13)), 0,  8) -- 11797
,( 9, E,0,0,((20,23),(18,21),( 2, 3),(20,23),(20,23),(12,15)), 0,  8) -- 11798
,( 9, E,0,0,((22,25),(20,23),( 4, 5),(22,25),(22,25),(14,17)), 0,  8) -- 11799
,( 9, E,0,0,((24,27),(22,25),( 6, 7),(24,27),(24,27),(16,19)), 0,  8) -- 11800
,( 9, E,0,0,((18,21),(16,19),( 0, 1),(18,21),(22,25),( 4, 7)), 0,  8) -- 11801
,( 9, E,0,0,((20,23),(18,21),( 2, 3),(20,23),(24,27),( 6, 9)), 0,  8) -- 11802
,( 9, E,0,0,((22,25),(20,23),( 4, 5),(22,25),(26,29),( 8,11)), 0,  8) -- 11803
,( 9, E,0,0,((24,27),(22,25),( 6, 7),(24,27),(28,31),(10,13)), 0,  8) -- 11804
,( 9, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 11805
,( 9, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 11806
,( 9, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 11807
,( 9, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 11808
,( 9, E,0,0,((14,17),(14,17),( 0, 1),(18,21),(20,23),(99,99)), 0,  8) -- 11809
,( 9, E,0,0,((16,19),(16,19),( 2, 3),(20,23),(22,25),(99,99)), 0,  8) -- 11810
,( 9, E,0,0,((18,21),(18,21),( 4, 5),(22,25),(24,27),(99,99)), 0,  8) -- 11811
,( 9, E,0,0,((20,23),(20,23),( 6, 7),(24,27),(26,29),(99,99)), 0,  8) -- 11812
,( 9, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(16,19),(99,99)), 0,  7) -- 11813
,( 9, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(18,21),(99,99)), 0,  7) -- 11814
,( 9, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(20,23),(99,99)), 0,  7) -- 11815
,( 9, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(22,25),(99,99)), 0,  7) -- 11816
,( 9, E,0,0,((14,17),(14,17),( 0, 1),(20,23),(24,27),(99,99)), 0,  7) -- 11817
,( 9, E,0,0,((16,19),(16,19),( 2, 3),(22,25),(26,29),(99,99)), 0,  7) -- 11818
,( 9, E,0,0,((18,21),(18,21),( 4, 5),(24,27),(28,31),(99,99)), 0,  7) -- 11819
,( 9, E,0,0,((20,23),(20,23),( 6, 7),(26,29),(30,33),(99,99)), 0,  7) -- 11820
,( 9, E,0,1,((10,13),(12,15),( 0, 1),(20,23),(99,99),(99,99)), 0,  7) -- 11821
,( 9, E,0,1,((12,15),(14,17),( 2, 3),(22,25),(99,99),(99,99)), 0,  7) -- 11822
,( 9, E,0,1,((14,17),(16,19),( 4, 5),(24,27),(99,99),(99,99)), 0,  7) -- 11823
,( 9, E,0,1,((16,19),(18,21),( 6, 7),(26,29),(99,99),(99,99)), 0,  7) -- 11824
,( 9, E,0,1,((16,19),(16,19),( 0, 1),(16,19),(99,99),(99,99)), 0,  7) -- 11825
,( 9, E,0,1,((18,21),(18,21),( 2, 3),(18,21),(99,99),(99,99)), 0,  7) -- 11826
,( 9, E,0,1,((20,23),(20,23),( 4, 5),(20,23),(99,99),(99,99)), 0,  7) -- 11827
,( 9, E,0,1,((22,25),(22,25),( 6, 7),(22,25),(99,99),(99,99)), 0,  7) -- 11828
,( 9, E,0,1,((12,15),(14,17),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 11829
,( 9, E,0,1,((14,17),(16,19),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 11830
,( 9, E,0,1,((16,19),(18,21),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 11831
,( 9, E,0,1,((18,21),(20,23),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 11832
,( 9, E,0,1,(( 8,11),(12,15),( 0, 1),(16,19),(99,99),(99,99)), 0,  6) -- 11833
,( 9, E,0,1,((10,13),(14,17),( 2, 3),(18,21),(99,99),(99,99)), 0,  6) -- 11834
,( 9, E,0,1,((12,15),(16,19),( 4, 5),(20,23),(99,99),(99,99)), 0,  6) -- 11835
,( 9, E,0,1,((14,17),(18,21),( 6, 7),(22,25),(99,99),(99,99)), 0,  6) -- 11836
,( 9, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 11837
,( 9, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 11838
,( 9, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 11839
,( 9, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 11840
,( 9, E,0,1,(( 6, 9),(10,13),( 0, 1),(20,23),(99,99),(99,99)), 0,  5) -- 11841
,( 9, E,0,1,(( 8,11),(12,15),( 2, 3),(22,25),(99,99),(99,99)), 0,  5) -- 11842
,( 9, E,0,1,((10,13),(14,17),( 4, 5),(24,27),(99,99),(99,99)), 0,  5) -- 11843
,( 9, E,0,1,((12,15),(16,19),( 6, 7),(26,29),(99,99),(99,99)), 0,  5) -- 11844
,( 9, E,0,1,((14,17),(16,19),( 0, 1),(14,15),(99,99),(99,99)), 0,  5) -- 11845
,( 9, E,0,1,((16,19),(18,21),( 2, 3),(16,17),(99,99),(99,99)), 0,  5) -- 11846
,( 9, E,0,1,((18,21),(20,23),( 4, 5),(18,19),(99,99),(99,99)), 0,  5) -- 11847
,( 9, E,0,1,((20,23),(22,25),( 6, 7),(20,21),(99,99),(99,99)), 0,  5) -- 11848
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 31) -- 11849
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 31) -- 11850
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 1, 31) -- 11851
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 1, 31) -- 11852
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 1, 31) -- 11853
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 1, 31) -- 11854
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 1, 31) -- 11855
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 1, 31) -- 11856
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 11857
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 11858
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 11859
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 11860
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 11861
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 11862
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 11863
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 11864
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 11865
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 11866
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 11867
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 11868
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 11869
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 11870
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 11871
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 11872
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 11873
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 11874
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 11875
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 11876
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 11877
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 11878
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 11879
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 11880
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 31) -- 11881
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 31) -- 11882
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 31) -- 11883
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 31) -- 11884
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 31) -- 11885
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 31) -- 11886
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 31) -- 11887
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 31) -- 11888
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 11889
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 11890
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 11891
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 11892
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 11893
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 11894
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 11895
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 11896
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 11897
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 11898
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 11899
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 11900
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 11901
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 11902
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 11903
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 11904
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 11905
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 11906
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 11907
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 11908
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 11909
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 11910
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 11911
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 11912
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 28) -- 11913
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 28) -- 11914
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 1, 28) -- 11915
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 1, 28) -- 11916
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 1, 28) -- 11917
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 1, 28) -- 11918
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 1, 28) -- 11919
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 1, 28) -- 11920
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(17,17),( 8, 8)), 1, 28) -- 11921
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(18,18),( 9, 9)), 1, 28) -- 11922
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(19,19),(10,10)), 1, 28) -- 11923
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(20,20),(11,11)), 1, 28) -- 11924
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(21,21),(12,12)), 1, 28) -- 11925
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(22,22),(13,13)), 1, 28) -- 11926
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(23,23),(14,14)), 1, 28) -- 11927
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(24,24),(15,15)), 1, 28) -- 11928
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 27) -- 11929
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 27) -- 11930
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 27) -- 11931
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(10,10)), 1, 27) -- 11932
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(11,11)), 1, 27) -- 11933
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(12,12)), 1, 27) -- 11934
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(13,13)), 1, 27) -- 11935
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(14,14)), 1, 27) -- 11936
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 26) -- 11937
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 26) -- 11938
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 26) -- 11939
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 26) -- 11940
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 26) -- 11941
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 26) -- 11942
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 26) -- 11943
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 26) -- 11944
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 25) -- 11945
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 25) -- 11946
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 25) -- 11947
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 25) -- 11948
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 25) -- 11949
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 25) -- 11950
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 25) -- 11951
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 25) -- 11952
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 25) -- 11953
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 25) -- 11954
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 25) -- 11955
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 25) -- 11956
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 25) -- 11957
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 25) -- 11958
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 25) -- 11959
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 25) -- 11960
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 24) -- 11961
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 24) -- 11962
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 24) -- 11963
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 24) -- 11964
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 24) -- 11965
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 24) -- 11966
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 24) -- 11967
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 24) -- 11968
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 24) -- 11969
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 24) -- 11970
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 24) -- 11971
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 24) -- 11972
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 24) -- 11973
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 24) -- 11974
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 24) -- 11975
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 24) -- 11976
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 23) -- 11977
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 23) -- 11978
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 23) -- 11979
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 23) -- 11980
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 23) -- 11981
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 23) -- 11982
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 23) -- 11983
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 23) -- 11984
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 23) -- 11985
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 23) -- 11986
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 23) -- 11987
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 23) -- 11988
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 23) -- 11989
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 23) -- 11990
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 23) -- 11991
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 23) -- 11992
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 22) -- 11993
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 22) -- 11994
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 22) -- 11995
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 22) -- 11996
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 22) -- 11997
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 22) -- 11998
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 22) -- 11999
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 22) -- 12000
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 22) -- 12001
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 22) -- 12002
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 22) -- 12003
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 22) -- 12004
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 22) -- 12005
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 22) -- 12006
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 22) -- 12007
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 22) -- 12008
,( 10, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 21) -- 12009
,( 10, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 21) -- 12010
,( 10, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 21) -- 12011
,( 10, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 21) -- 12012
,( 10, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 21) -- 12013
,( 10, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 21) -- 12014
,( 10, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 21) -- 12015
,( 10, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 21) -- 12016
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(16,16),( 6, 6)), 1, 21) -- 12017
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(17,17),( 7, 7)), 1, 21) -- 12018
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(18,18),( 8, 8)), 1, 21) -- 12019
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(19,19),( 9, 9)), 1, 21) -- 12020
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(20,20),(10,10)), 1, 21) -- 12021
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(21,21),(11,11)), 1, 21) -- 12022
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(22,22),(12,12)), 1, 21) -- 12023
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(23,23),(13,13)), 1, 21) -- 12024
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 20) -- 12025
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 20) -- 12026
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 20) -- 12027
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 20) -- 12028
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 20) -- 12029
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 20) -- 12030
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 20) -- 12031
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 20) -- 12032
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 20) -- 12033
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 20) -- 12034
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 20) -- 12035
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 20) -- 12036
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 20) -- 12037
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 20) -- 12038
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 20) -- 12039
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 20) -- 12040
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 19) -- 12041
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 19) -- 12042
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 19) -- 12043
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(19,19),(10,10)), 1, 19) -- 12044
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(20,20),(11,11)), 1, 19) -- 12045
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(21,21),(12,12)), 1, 19) -- 12046
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(22,22),(13,13)), 1, 19) -- 12047
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(23,23),(14,14)), 1, 19) -- 12048
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 12049
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 12050
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 12051
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 12052
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 12053
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 12054
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 12055
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 12056
,( 10, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 19) -- 12057
,( 10, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 19) -- 12058
,( 10, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 19) -- 12059
,( 10, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 19) -- 12060
,( 10, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 19) -- 12061
,( 10, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 19) -- 12062
,( 10, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 19) -- 12063
,( 10, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 19) -- 12064
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(16,16),( 6, 6)), 1, 19) -- 12065
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(17,17),( 7, 7)), 1, 19) -- 12066
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(18,18),( 8, 8)), 1, 19) -- 12067
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(19,19),( 9, 9)), 1, 19) -- 12068
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(20,20),(10,10)), 1, 19) -- 12069
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(21,21),(11,11)), 1, 19) -- 12070
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(22,22),(12,12)), 1, 19) -- 12071
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(23,23),(13,13)), 1, 19) -- 12072
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 18) -- 12073
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 18) -- 12074
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 18) -- 12075
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 18) -- 12076
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 18) -- 12077
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 18) -- 12078
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 18) -- 12079
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 18) -- 12080
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 18) -- 12081
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 18) -- 12082
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 18) -- 12083
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 18) -- 12084
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 18) -- 12085
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(10,10)), 1, 18) -- 12086
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(11,11)), 1, 18) -- 12087
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(12,12)), 1, 18) -- 12088
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 12089
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 12090
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 12091
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 12092
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 12093
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 12094
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 12095
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 12096
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 12097
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 12098
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 12099
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 12100
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 12101
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 12102
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 12103
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 12104
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 17) -- 12105
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 17) -- 12106
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 17) -- 12107
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 17) -- 12108
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 17) -- 12109
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 17) -- 12110
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 17) -- 12111
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 17) -- 12112
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 12113
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 12114
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 12115
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 12116
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 12117
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 12118
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 12119
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 12120
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 12121
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 12122
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 12123
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 12124
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 12125
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 12126
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 12127
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 12128
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 17) -- 12129
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 17) -- 12130
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 17) -- 12131
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 17) -- 12132
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 17) -- 12133
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(10,10)), 1, 17) -- 12134
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(11,11)), 1, 17) -- 12135
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(12,12)), 1, 17) -- 12136
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 12137
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 12138
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 12139
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 12140
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 12141
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 12142
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 12143
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 12144
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(15,15),( 5, 5)), 1, 16) -- 12145
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(16,16),( 6, 6)), 1, 16) -- 12146
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(17,17),( 7, 7)), 1, 16) -- 12147
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(18,18),( 8, 8)), 1, 16) -- 12148
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(19,19),( 9, 9)), 1, 16) -- 12149
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(20,20),(10,10)), 1, 16) -- 12150
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(21,21),(11,11)), 1, 16) -- 12151
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(22,22),(12,12)), 1, 16) -- 12152
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 12153
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 12154
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 12155
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 12156
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 12157
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 12158
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 12159
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 12160
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 16) -- 12161
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 16) -- 12162
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 16) -- 12163
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 16) -- 12164
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 16) -- 12165
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 16) -- 12166
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 16) -- 12167
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 16) -- 12168
,( 10, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 16) -- 12169
,( 10, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 16) -- 12170
,( 10, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 16) -- 12171
,( 10, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 16) -- 12172
,( 10, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 16) -- 12173
,( 10, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 16) -- 12174
,( 10, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(10,10)), 1, 16) -- 12175
,( 10, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(11,11)), 1, 16) -- 12176
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 12177
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 12178
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 12179
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 12180
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 12181
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 12182
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 12183
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 12184
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 16) -- 12185
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 16) -- 12186
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 16) -- 12187
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 16) -- 12188
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 16) -- 12189
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 16) -- 12190
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 16) -- 12191
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 16) -- 12192
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 15) -- 12193
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 15) -- 12194
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 15) -- 12195
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 15) -- 12196
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 15) -- 12197
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 15) -- 12198
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(10,10)), 1, 15) -- 12199
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(11,11)), 1, 15) -- 12200
,( 10, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 12201
,( 10, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 12202
,( 10, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 12203
,( 10, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 12204
,( 10, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 12205
,( 10, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 12206
,( 10, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 12207
,( 10, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 12208
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 4, 4)), 1, 15) -- 12209
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 5, 5)), 1, 15) -- 12210
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 6, 6)), 1, 15) -- 12211
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 7, 7)), 1, 15) -- 12212
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 8, 8)), 1, 15) -- 12213
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),( 9, 9)), 1, 15) -- 12214
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(10,10)), 1, 15) -- 12215
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(11,11)), 1, 15) -- 12216
,( 10, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 15) -- 12217
,( 10, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 15) -- 12218
,( 10, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 15) -- 12219
,( 10, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 15) -- 12220
,( 10, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 15) -- 12221
,( 10, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 15) -- 12222
,( 10, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 15) -- 12223
,( 10, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 15) -- 12224
,( 10, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(14,14),( 4, 4)), 1, 15) -- 12225
,( 10, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(15,15),( 5, 5)), 1, 15) -- 12226
,( 10, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(16,16),( 6, 6)), 1, 15) -- 12227
,( 10, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(17,17),( 7, 7)), 1, 15) -- 12228
,( 10, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(18,18),( 8, 8)), 1, 15) -- 12229
,( 10, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(19,19),( 9, 9)), 1, 15) -- 12230
,( 10, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(20,20),(10,10)), 1, 15) -- 12231
,( 10, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(21,21),(11,11)), 1, 15) -- 12232
,( 10, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 12233
,( 10, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 12234
,( 10, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 12235
,( 10, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 12236
,( 10, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 12237
,( 10, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 12238
,( 10, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 12239
,( 10, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 12240
,( 10, E,0,0,((36,37),(27,27),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 14) -- 12241
,( 10, E,0,0,((38,39),(29,29),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 14) -- 12242
,( 10, E,0,0,((40,41),(31,31),( 5, 5),(20,20),(18,19),( 8,11)), 1, 14) -- 12243
,( 10, E,0,0,((42,43),(33,33),( 7, 7),(22,22),(20,21),(10,13)), 1, 14) -- 12244
,( 10, E,0,0,((36,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 13) -- 12245
,( 10, E,0,0,((38,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 13) -- 12246
,( 10, E,0,0,((40,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 13) -- 12247
,( 10, E,0,0,((42,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 13) -- 12248
,( 10, E,0,0,((38,38),(27,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 13) -- 12249
,( 10, E,0,0,((40,40),(29,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 13) -- 12250
,( 10, E,0,0,((42,42),(31,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 13) -- 12251
,( 10, E,0,0,((44,44),(33,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 13) -- 12252
,( 10, E,0,0,((36,39),(27,27),( 1, 1),(16,16),(16,16),( 6, 9)), 1, 13) -- 12253
,( 10, E,0,0,((38,41),(29,29),( 3, 3),(18,18),(18,18),( 8,11)), 1, 13) -- 12254
,( 10, E,0,0,((40,43),(31,31),( 5, 5),(20,20),(20,20),(10,13)), 1, 13) -- 12255
,( 10, E,0,0,((42,45),(33,33),( 7, 7),(22,22),(22,22),(12,15)), 1, 13) -- 12256
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 12) -- 12257
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 12) -- 12258
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),( 8,11)), 1, 12) -- 12259
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(10,13)), 1, 12) -- 12260
,( 10, E,0,0,((38,39),(27,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 12261
,( 10, E,0,0,((40,41),(29,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 12262
,( 10, E,0,0,((42,43),(31,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 12263
,( 10, E,0,0,((44,45),(33,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 12264
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 12265
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 12266
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 12267
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 12268
,( 10, E,0,0,((36,39),(26,27),( 0, 0),(13,13),(12,13),( 2, 5)), 1, 11) -- 12269
,( 10, E,0,0,((38,41),(28,29),( 2, 2),(15,15),(14,15),( 4, 7)), 1, 11) -- 12270
,( 10, E,0,0,((40,43),(30,31),( 4, 4),(17,17),(16,17),( 6, 9)), 1, 11) -- 12271
,( 10, E,0,0,((42,45),(32,33),( 6, 6),(19,19),(18,19),( 8,11)), 1, 11) -- 12272
,( 10, E,0,0,((38,39),(27,27),( 0, 0),(13,13),(11,11),( 0, 3)), 1, 11) -- 12273
,( 10, E,0,0,((40,41),(29,29),( 2, 2),(15,15),(13,13),( 2, 5)), 1, 11) -- 12274
,( 10, E,0,0,((42,43),(31,31),( 4, 4),(17,17),(15,15),( 4, 7)), 1, 11) -- 12275
,( 10, E,0,0,((44,45),(33,33),( 6, 6),(19,19),(17,17),( 6, 9)), 1, 11) -- 12276
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(13,13),(10,11),( 0, 3)), 1, 11) -- 12277
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(15,15),(12,13),( 2, 5)), 1, 11) -- 12278
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(17,17),(14,15),( 4, 7)), 1, 11) -- 12279
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(19,19),(16,17),( 6, 9)), 1, 11) -- 12280
,( 10, E,0,0,((38,41),(28,28),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 11) -- 12281
,( 10, E,0,0,((40,43),(30,30),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 11) -- 12282
,( 10, E,0,0,((42,45),(32,32),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 11) -- 12283
,( 10, E,0,0,((44,47),(34,34),( 6, 6),(19,19),(18,18),( 8,11)), 1, 11) -- 12284
,( 10, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(14,15),( 8,11)), 1, 11) -- 12285
,( 10, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(16,17),(10,13)), 1, 11) -- 12286
,( 10, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(18,19),(12,15)), 1, 11) -- 12287
,( 10, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(20,21),(14,17)), 1, 11) -- 12288
,( 10, E,0,0,((36,39),(26,27),( 0, 0),(14,14),(13,13),( 6, 7)), 1, 11) -- 12289
,( 10, E,0,0,((38,41),(28,29),( 2, 2),(16,16),(15,15),( 8, 9)), 1, 11) -- 12290
,( 10, E,0,0,((40,43),(30,31),( 4, 4),(18,18),(17,17),(10,11)), 1, 11) -- 12291
,( 10, E,0,0,((42,45),(32,33),( 6, 6),(20,20),(19,19),(12,13)), 1, 11) -- 12292
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 12293
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 12294
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 10) -- 12295
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 10) -- 12296
,( 10, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 10) -- 12297
,( 10, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 10) -- 12298
,( 10, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 10) -- 12299
,( 10, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(18,19),( 8,11)), 1, 10) -- 12300
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 8,11)), 1, 10) -- 12301
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(10,13)), 1, 10) -- 12302
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(12,15)), 1, 10) -- 12303
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(14,17)), 1, 10) -- 12304
,( 10, E,0,0,((40,43),(28,29),( 0, 1),(12,13),(10,11),( 2, 5)), 1, 10) -- 12305
,( 10, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(12,13),( 4, 7)), 1, 10) -- 12306
,( 10, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(14,15),( 6, 9)), 1, 10) -- 12307
,( 10, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(16,17),( 8,11)), 1, 10) -- 12308
,( 10, E,0,0,((38,41),(28,29),( 0, 1),(13,13),(12,13),( 4, 7)), 1, 10) -- 12309
,( 10, E,0,0,((40,43),(30,31),( 2, 3),(15,15),(14,15),( 6, 9)), 1, 10) -- 12310
,( 10, E,0,0,((42,45),(32,33),( 4, 5),(17,17),(16,17),( 8,11)), 1, 10) -- 12311
,( 10, E,0,0,((44,47),(34,35),( 6, 7),(19,19),(18,19),(10,13)), 1, 10) -- 12312
,( 10, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(11,11),( 0, 3)), 1, 10) -- 12313
,( 10, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(13,13),( 2, 5)), 1, 10) -- 12314
,( 10, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(15,15),( 4, 7)), 1, 10) -- 12315
,( 10, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(17,17),( 6, 9)), 1, 10) -- 12316
,( 10, E,0,0,((42,43),(30,30),( 1, 1),(14,14),(10,11),( 0, 3)), 1, 10) -- 12317
,( 10, E,0,0,((44,45),(32,32),( 3, 3),(16,16),(12,13),( 2, 5)), 1, 10) -- 12318
,( 10, E,0,0,((46,47),(34,34),( 5, 5),(18,18),(14,15),( 4, 7)), 1, 10) -- 12319
,( 10, E,0,0,((48,49),(36,36),( 7, 7),(20,20),(16,17),( 6, 9)), 1, 10) -- 12320
,( 10, E,0,0,((42,42),(29,29),( 1, 1),(14,14),(12,13),( 4, 7)), 1, 10) -- 12321
,( 10, E,0,0,((44,44),(31,31),( 3, 3),(16,16),(14,15),( 6, 9)), 1, 10) -- 12322
,( 10, E,0,0,((46,46),(33,33),( 5, 5),(18,18),(16,17),( 8,11)), 1, 10) -- 12323
,( 10, E,0,0,((48,48),(35,35),( 7, 7),(20,20),(18,19),(10,13)), 1, 10) -- 12324
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),( 6, 9)), 1,  9) -- 12325
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),( 8,11)), 1,  9) -- 12326
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(10,13)), 1,  9) -- 12327
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(12,15)), 1,  9) -- 12328
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 2, 5)), 1,  9) -- 12329
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 4, 7)), 1,  9) -- 12330
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 6, 9)), 1,  9) -- 12331
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 8,11)), 1,  9) -- 12332
,( 10, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(12,13),( 8,11)), 1,  9) -- 12333
,( 10, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(14,15),(10,13)), 1,  9) -- 12334
,( 10, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(16,17),(12,15)), 1,  9) -- 12335
,( 10, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(18,19),(14,17)), 1,  9) -- 12336
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(12,13),( 6, 9)), 1,  9) -- 12337
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(14,15),( 8,11)), 1,  9) -- 12338
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(16,17),(10,13)), 1,  9) -- 12339
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(18,19),(12,15)), 1,  9) -- 12340
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(14,15),( 8,11)), 1,  9) -- 12341
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(16,17),(10,13)), 1,  9) -- 12342
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(18,19),(12,15)), 1,  9) -- 12343
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(20,21),(14,17)), 1,  9) -- 12344
,( 10, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 6, 9)), 1,  9) -- 12345
,( 10, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 8,11)), 1,  9) -- 12346
,( 10, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),(10,13)), 1,  9) -- 12347
,( 10, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),(12,15)), 1,  9) -- 12348
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 12349
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 12350
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 12351
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 12352
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 6, 9)), 1,  9) -- 12353
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 8,11)), 1,  9) -- 12354
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(10,13)), 1,  9) -- 12355
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(12,15)), 1,  9) -- 12356
,( 10, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1,  9) -- 12357
,( 10, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1,  9) -- 12358
,( 10, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1,  9) -- 12359
,( 10, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1,  9) -- 12360
,( 10, E,0,0,((40,43),(28,29),( 0, 1),(14,14),(12,13),( 8,11)), 1,  9) -- 12361
,( 10, E,0,0,((42,45),(30,31),( 2, 3),(16,16),(14,15),(10,13)), 1,  9) -- 12362
,( 10, E,0,0,((44,47),(32,33),( 4, 5),(18,18),(16,17),(12,15)), 1,  9) -- 12363
,( 10, E,0,0,((46,49),(34,35),( 6, 7),(20,20),(18,19),(14,17)), 1,  9) -- 12364
,( 10, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(12,13),(10,13)), 1,  9) -- 12365
,( 10, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(14,15),(12,15)), 1,  9) -- 12366
,( 10, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(16,17),(14,17)), 1,  9) -- 12367
,( 10, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(18,19),(16,19)), 1,  9) -- 12368
,( 10, E,0,0,((40,43),(29,29),( 0, 0),(12,12),( 8, 9),( 0, 3)), 1,  9) -- 12369
,( 10, E,0,0,((42,45),(31,31),( 2, 2),(14,14),(10,11),( 2, 5)), 1,  9) -- 12370
,( 10, E,0,0,((44,47),(33,33),( 4, 4),(16,16),(12,13),( 4, 7)), 1,  9) -- 12371
,( 10, E,0,0,((46,49),(35,35),( 6, 6),(18,18),(14,15),( 6, 9)), 1,  9) -- 12372
,( 10, E,0,0,((42,43),(29,29),( 0, 1),(13,13),(12,12),( 4, 7)), 1,  9) -- 12373
,( 10, E,0,0,((44,45),(31,31),( 2, 3),(15,15),(14,14),( 6, 9)), 1,  9) -- 12374
,( 10, E,0,0,((46,47),(33,33),( 4, 5),(17,17),(16,16),( 8,11)), 1,  9) -- 12375
,( 10, E,0,0,((48,49),(35,35),( 6, 7),(19,19),(18,18),(10,13)), 1,  9) -- 12376
,( 10, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 2, 5)), 1,  9) -- 12377
,( 10, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 4, 7)), 1,  9) -- 12378
,( 10, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 6, 9)), 1,  9) -- 12379
,( 10, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),( 8,11)), 1,  9) -- 12380
,( 10, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(14,15),(14,17)), 1,  9) -- 12381
,( 10, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(16,17),(16,19)), 1,  9) -- 12382
,( 10, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(18,19),(18,21)), 1,  9) -- 12383
,( 10, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(20,21),(20,23)), 1,  9) -- 12384
,( 10, E,0,0,((44,47),(32,32),( 1, 1),(13,13),(10,11),( 2, 5)), 1,  9) -- 12385
,( 10, E,0,0,((46,49),(34,34),( 3, 3),(15,15),(12,13),( 4, 7)), 1,  9) -- 12386
,( 10, E,0,0,((48,51),(36,36),( 5, 5),(17,17),(14,15),( 6, 9)), 1,  9) -- 12387
,( 10, E,0,0,((50,53),(38,38),( 7, 7),(19,19),(16,17),( 8,11)), 1,  9) -- 12388
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(14,14),(12,13),( 2, 5)), 1,  9) -- 12389
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(16,16),(14,15),( 4, 7)), 1,  9) -- 12390
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(18,18),(16,17),( 6, 9)), 1,  9) -- 12391
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(20,20),(18,19),( 8,11)), 1,  9) -- 12392
,( 10, E,0,0,((42,43),(30,30),( 1, 1),(14,15),(14,15),(12,15)), 1,  9) -- 12393
,( 10, E,0,0,((44,45),(32,32),( 3, 3),(16,17),(16,17),(14,17)), 1,  9) -- 12394
,( 10, E,0,0,((46,47),(34,34),( 5, 5),(18,19),(18,19),(16,19)), 1,  9) -- 12395
,( 10, E,0,0,((48,49),(36,36),( 7, 7),(20,21),(20,21),(18,21)), 1,  9) -- 12396
,( 10, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(16,17),(16,16)), 1,  9) -- 12397
,( 10, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(18,19),(18,18)), 1,  9) -- 12398
,( 10, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(20,21),(20,20)), 1,  9) -- 12399
,( 10, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(22,23),(22,22)), 1,  9) -- 12400
,( 10, E,0,0,((46,46),(31,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 12401
,( 10, E,0,0,((48,48),(33,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 12402
,( 10, E,0,0,((50,50),(35,35),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 12403
,( 10, E,0,0,((52,52),(37,37),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 12404
,( 10, E,0,0,((42,45),(30,31),( 0, 1),(13,13),(12,12),( 2, 5)), 1,  9) -- 12405
,( 10, E,0,0,((44,47),(32,33),( 2, 3),(15,15),(14,14),( 4, 7)), 1,  9) -- 12406
,( 10, E,0,0,((46,49),(34,35),( 4, 5),(17,17),(16,16),( 6, 9)), 1,  9) -- 12407
,( 10, E,0,0,((48,51),(36,37),( 6, 7),(19,19),(18,18),( 8,11)), 1,  9) -- 12408
,( 10, E,0,0,((42,42),(29,29),( 0, 0),(14,14),(12,12),( 2, 5)), 1,  9) -- 12409
,( 10, E,0,0,((44,44),(31,31),( 2, 2),(16,16),(14,14),( 4, 7)), 1,  9) -- 12410
,( 10, E,0,0,((46,46),(33,33),( 4, 4),(18,18),(16,16),( 6, 9)), 1,  9) -- 12411
,( 10, E,0,0,((48,48),(35,35),( 6, 6),(20,20),(18,18),( 8,11)), 1,  9) -- 12412
,( 10, E,0,0,((42,45),(30,30),( 0, 1),(12,13),(10,11),( 0, 1)), 1,  9) -- 12413
,( 10, E,0,0,((44,47),(32,32),( 2, 3),(14,15),(12,13),( 2, 3)), 1,  9) -- 12414
,( 10, E,0,0,((46,49),(34,34),( 4, 5),(16,17),(14,15),( 4, 5)), 1,  9) -- 12415
,( 10, E,0,0,((48,51),(36,36),( 6, 7),(18,19),(16,17),( 6, 7)), 1,  9) -- 12416
,( 10, E,0,0,((40,43),(28,29),( 0, 0),(12,13),(10,11),( 0, 1)), 1,  9) -- 12417
,( 10, E,0,0,((42,45),(30,31),( 2, 2),(14,15),(12,13),( 2, 3)), 1,  9) -- 12418
,( 10, E,0,0,((44,47),(32,33),( 4, 4),(16,17),(14,15),( 4, 5)), 1,  9) -- 12419
,( 10, E,0,0,((46,49),(34,35),( 6, 6),(18,19),(16,17),( 6, 7)), 1,  9) -- 12420
,( 10, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(12,15),(11,11)), 1,  8) -- 12421
,( 10, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(14,17),(13,13)), 1,  8) -- 12422
,( 10, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(16,19),(15,15)), 1,  8) -- 12423
,( 10, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(18,21),(17,17)), 1,  8) -- 12424
,( 10, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(18,21)), 1,  8) -- 12425
,( 10, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(20,23)), 1,  8) -- 12426
,( 10, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(22,23)), 1,  8) -- 12427
,( 10, E,0,0,((46,49),(30,33),( 0, 1),(10,13),( 8,11),(99,99)), 1,  8) -- 12428
,( 10, E,0,0,((48,51),(32,35),( 2, 3),(12,15),(10,13),(99,99)), 1,  8) -- 12429
,( 10, E,0,0,((50,53),(34,37),( 4, 5),(14,17),(12,15),(99,99)), 1,  8) -- 12430
,( 10, E,0,0,((52,55),(36,39),( 6, 7),(16,19),(14,17),(99,99)), 1,  8) -- 12431
,( 10, E,0,0,((48,51),(32,35),( 0, 1),(12,15),(12,15),(99,99)), 1,  7) -- 12432
,( 10, E,0,0,((50,53),(34,37),( 2, 3),(14,17),(14,17),(99,99)), 1,  7) -- 12433
,( 10, E,0,0,((52,55),(36,39),( 4, 5),(16,19),(16,19),(99,99)), 1,  7) -- 12434
,( 10, E,0,0,((54,57),(38,41),( 6, 7),(18,21),(18,21),(99,99)), 1,  7) -- 12435
,( 10, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(16,19),(99,99)), 1,  7) -- 12436
,( 10, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(18,21),(99,99)), 1,  7) -- 12437
,( 10, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(20,23),(99,99)), 1,  7) -- 12438
,( 10, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(22,25),(99,99)), 1,  7) -- 12439
,( 10, E,0,1,((48,51),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  7) -- 12440
,( 10, E,0,1,((50,53),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  7) -- 12441
,( 10, E,0,1,((52,55),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  7) -- 12442
,( 10, E,0,1,((54,57),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  7) -- 12443
,( 10, E,0,1,((44,47),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 12444
,( 10, E,0,1,((46,49),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 12445
,( 10, E,0,1,((48,51),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 12446
,( 10, E,0,1,((50,53),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 12447
,( 10, E,0,1,((50,53),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  6) -- 12448
,( 10, E,0,1,((52,55),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  6) -- 12449
,( 10, E,0,1,((54,57),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  6) -- 12450
,( 10, E,0,1,((56,59),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  6) -- 12451
,( 10, E,0,1,((48,51),(30,33),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 12452
,( 10, E,0,1,((50,53),(32,35),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 12453
,( 10, E,0,1,((52,55),(34,37),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 12454
,( 10, E,0,1,((54,57),(36,39),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 12455
,( 10, E,0,1,((52,55),(32,35),( 0, 1),(14,17),(99,99),(99,99)), 1,  6) -- 12456
,( 10, E,0,1,((54,57),(34,37),( 2, 3),(16,19),(99,99),(99,99)), 1,  6) -- 12457
,( 10, E,0,1,((56,59),(36,39),( 4, 5),(18,21),(99,99),(99,99)), 1,  6) -- 12458
,( 10, E,0,1,((58,61),(38,41),( 6, 7),(20,23),(99,99),(99,99)), 1,  6) -- 12459
,( 10, E,0,1,((36,39),(26,27),( 0, 1),(18,19),(99,99),(99,99)), 1,  5) -- 12460
,( 10, E,0,1,((38,41),(28,29),( 2, 3),(20,21),(99,99),(99,99)), 1,  5) -- 12461
,( 10, E,0,1,((40,43),(30,31),( 4, 5),(22,23),(99,99),(99,99)), 1,  5) -- 12462
,( 10, E,0,1,((42,45),(32,33),( 6, 7),(24,25),(99,99),(99,99)), 1,  5) -- 12463
,( 10, E,0,1,((46,49),(30,33),( 1, 1),(18,18),(99,99),(99,99)), 1,  5) -- 12464
,( 10, E,0,1,((48,51),(32,35),( 3, 3),(20,20),(99,99),(99,99)), 1,  5) -- 12465
,( 10, E,0,1,((50,53),(34,37),( 5, 5),(22,22),(99,99),(99,99)), 1,  5) -- 12466
,( 10, E,0,1,((52,55),(36,39),( 7, 7),(24,24),(99,99),(99,99)), 1,  5) -- 12467
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 12468
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 12469
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 12470
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 12471
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 12472
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 12473
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 12474
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 12475
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 12476
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 12477
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 12478
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 12479
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 12480
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 12481
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 12482
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 12483
,( 10, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 12484
,( 10, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 12485
,( 10, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 12486
,( 10, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 12487
,( 10, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 12488
,( 10, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 12489
,( 10, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 12490
,( 10, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 12491
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 31) -- 12492
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 31) -- 12493
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(10,10)), 0, 31) -- 12494
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(11,11)), 0, 31) -- 12495
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(12,12)), 0, 31) -- 12496
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(13,13)), 0, 31) -- 12497
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(14,14)), 0, 31) -- 12498
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(15,15)), 0, 31) -- 12499
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 12500
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 12501
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 12502
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 12503
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 12504
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 12505
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 12506
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 12507
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 7, 7)), 0, 31) -- 12508
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 8, 8)), 0, 31) -- 12509
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),( 9, 9)), 0, 31) -- 12510
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(10,10)), 0, 31) -- 12511
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(11,11)), 0, 31) -- 12512
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(12,12)), 0, 31) -- 12513
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(13,13)), 0, 31) -- 12514
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(14,14)), 0, 31) -- 12515
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(17,17),( 8, 8)), 0, 31) -- 12516
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(18,18),( 9, 9)), 0, 31) -- 12517
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(19,19),(10,10)), 0, 31) -- 12518
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(20,20),(11,11)), 0, 31) -- 12519
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(21,21),(12,12)), 0, 31) -- 12520
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(22,22),(13,13)), 0, 31) -- 12521
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(23,23),(14,14)), 0, 31) -- 12522
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(24,24),(15,15)), 0, 31) -- 12523
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 12524
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 12525
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 12526
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 12527
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 12528
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 12529
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 12530
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 12531
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 30) -- 12532
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 30) -- 12533
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 30) -- 12534
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 30) -- 12535
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 30) -- 12536
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 30) -- 12537
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 30) -- 12538
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 30) -- 12539
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 29) -- 12540
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 29) -- 12541
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 29) -- 12542
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 29) -- 12543
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 29) -- 12544
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 29) -- 12545
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 29) -- 12546
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 29) -- 12547
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 27) -- 12548
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 27) -- 12549
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 27) -- 12550
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 27) -- 12551
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 27) -- 12552
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 27) -- 12553
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 27) -- 12554
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 27) -- 12555
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(17,17),( 9, 9)), 0, 25) -- 12556
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(18,18),(10,10)), 0, 25) -- 12557
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(19,19),(11,11)), 0, 25) -- 12558
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(20,20),(12,12)), 0, 25) -- 12559
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(21,21),(13,13)), 0, 25) -- 12560
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(22,22),(14,14)), 0, 25) -- 12561
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(23,23),(15,15)), 0, 25) -- 12562
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(24,24),(16,16)), 0, 25) -- 12563
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(17,17),( 8, 8)), 0, 24) -- 12564
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(18,18),( 9, 9)), 0, 24) -- 12565
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(19,19),(10,10)), 0, 24) -- 12566
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(20,20),(11,11)), 0, 24) -- 12567
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(21,21),(12,12)), 0, 24) -- 12568
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(22,22),(13,13)), 0, 24) -- 12569
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(23,23),(14,14)), 0, 24) -- 12570
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(24,24),(15,15)), 0, 24) -- 12571
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 24) -- 12572
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(10,10)), 0, 24) -- 12573
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(11,11)), 0, 24) -- 12574
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(12,12)), 0, 24) -- 12575
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(13,13)), 0, 24) -- 12576
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(14,14)), 0, 24) -- 12577
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(15,15)), 0, 24) -- 12578
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(16,16)), 0, 24) -- 12579
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 8, 8)), 0, 24) -- 12580
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),( 9, 9)), 0, 24) -- 12581
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(10,10)), 0, 24) -- 12582
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(11,11)), 0, 24) -- 12583
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(12,12)), 0, 24) -- 12584
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(13,13)), 0, 24) -- 12585
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(14,14)), 0, 24) -- 12586
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(15,15)), 0, 24) -- 12587
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(18,18),(10,10)), 0, 24) -- 12588
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(19,19),(11,11)), 0, 24) -- 12589
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(20,20),(12,12)), 0, 24) -- 12590
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(21,21),(13,13)), 0, 24) -- 12591
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(22,22),(14,14)), 0, 24) -- 12592
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(23,23),(15,15)), 0, 24) -- 12593
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(24,24),(16,16)), 0, 24) -- 12594
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(25,25),(17,17)), 0, 24) -- 12595
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 23) -- 12596
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 23) -- 12597
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 23) -- 12598
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 23) -- 12599
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 23) -- 12600
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 23) -- 12601
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 23) -- 12602
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 23) -- 12603
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(17,17),( 9, 9)), 0, 22) -- 12604
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(18,18),(10,10)), 0, 22) -- 12605
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(19,19),(11,11)), 0, 22) -- 12606
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(20,20),(12,12)), 0, 22) -- 12607
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(21,21),(13,13)), 0, 22) -- 12608
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(22,22),(14,14)), 0, 22) -- 12609
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(23,23),(15,15)), 0, 22) -- 12610
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(24,24),(16,16)), 0, 22) -- 12611
,( 10, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 22) -- 12612
,( 10, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 22) -- 12613
,( 10, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 22) -- 12614
,( 10, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 22) -- 12615
,( 10, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 22) -- 12616
,( 10, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 22) -- 12617
,( 10, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 22) -- 12618
,( 10, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 22) -- 12619
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 21) -- 12620
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 21) -- 12621
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 21) -- 12622
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 21) -- 12623
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 21) -- 12624
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 21) -- 12625
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 21) -- 12626
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 21) -- 12627
,( 10, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 21) -- 12628
,( 10, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 21) -- 12629
,( 10, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 21) -- 12630
,( 10, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 21) -- 12631
,( 10, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 21) -- 12632
,( 10, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 21) -- 12633
,( 10, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 21) -- 12634
,( 10, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 21) -- 12635
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 20) -- 12636
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 20) -- 12637
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 20) -- 12638
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 20) -- 12639
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 20) -- 12640
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 20) -- 12641
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 20) -- 12642
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 20) -- 12643
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 20) -- 12644
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 20) -- 12645
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 20) -- 12646
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 20) -- 12647
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 20) -- 12648
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 20) -- 12649
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 20) -- 12650
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 20) -- 12651
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 20) -- 12652
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 20) -- 12653
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 20) -- 12654
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 20) -- 12655
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 20) -- 12656
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 20) -- 12657
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 20) -- 12658
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 20) -- 12659
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 12660
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 12661
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 12662
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 12663
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 12664
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 12665
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 12666
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 12667
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 12668
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 12669
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 12670
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 12671
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 12672
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 12673
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 12674
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 12675
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 12676
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 12677
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 12678
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 12679
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 12680
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 12681
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 12682
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 12683
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 19) -- 12684
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 19) -- 12685
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 19) -- 12686
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 19) -- 12687
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 19) -- 12688
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 19) -- 12689
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 19) -- 12690
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 19) -- 12691
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 12692
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 12693
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 12694
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 12695
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 12696
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 12697
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 12698
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 12699
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 12700
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 12701
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 12702
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 12703
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 12704
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 12705
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 12706
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 12707
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 18) -- 12708
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(10,10)), 0, 18) -- 12709
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(11,11)), 0, 18) -- 12710
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(12,12)), 0, 18) -- 12711
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(13,13)), 0, 18) -- 12712
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(14,14)), 0, 18) -- 12713
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(15,15)), 0, 18) -- 12714
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(16,16)), 0, 18) -- 12715
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 12716
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 12717
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 12718
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 12719
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 12720
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 12721
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 12722
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 12723
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 18) -- 12724
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 18) -- 12725
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 18) -- 12726
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 18) -- 12727
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 18) -- 12728
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 18) -- 12729
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 18) -- 12730
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 18) -- 12731
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 12732
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 12733
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 12734
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 12735
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 12736
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 12737
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 12738
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 12739
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 12740
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 12741
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 12742
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 12743
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 12744
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 12745
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 12746
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 12747
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 17) -- 12748
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 17) -- 12749
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 17) -- 12750
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 17) -- 12751
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 17) -- 12752
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 17) -- 12753
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 17) -- 12754
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 17) -- 12755
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 12756
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 12757
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 12758
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 12759
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 12760
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 12761
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 12762
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 12763
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 17) -- 12764
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 17) -- 12765
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 17) -- 12766
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 17) -- 12767
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 17) -- 12768
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 17) -- 12769
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 17) -- 12770
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 17) -- 12771
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 17) -- 12772
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(10,10)), 0, 17) -- 12773
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(11,11)), 0, 17) -- 12774
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(12,12)), 0, 17) -- 12775
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(13,13)), 0, 17) -- 12776
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(14,14)), 0, 17) -- 12777
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(15,15)), 0, 17) -- 12778
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(16,16)), 0, 17) -- 12779
,( 10, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),( 9, 9)), 0, 17) -- 12780
,( 10, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(10,10)), 0, 17) -- 12781
,( 10, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(11,11)), 0, 17) -- 12782
,( 10, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(12,12)), 0, 17) -- 12783
,( 10, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(13,13)), 0, 17) -- 12784
,( 10, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(14,14)), 0, 17) -- 12785
,( 10, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(15,15)), 0, 17) -- 12786
,( 10, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(16,16)), 0, 17) -- 12787
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 12788
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 12789
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 12790
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 12791
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 12792
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 12793
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 12794
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 12795
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 12796
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 12797
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 12798
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 12799
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 12800
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 12801
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 12802
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 12803
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 16) -- 12804
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 16) -- 12805
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 16) -- 12806
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 16) -- 12807
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 16) -- 12808
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 16) -- 12809
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 16) -- 12810
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 16) -- 12811
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(10,10)), 0, 16) -- 12812
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(11,11)), 0, 16) -- 12813
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(12,12)), 0, 16) -- 12814
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(13,13)), 0, 16) -- 12815
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(14,14)), 0, 16) -- 12816
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(15,15)), 0, 16) -- 12817
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(16,16)), 0, 16) -- 12818
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(17,17)), 0, 16) -- 12819
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 12820
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 12821
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 12822
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 12823
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 12824
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 12825
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 12826
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 12827
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(10,10)), 0, 16) -- 12828
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(11,11)), 0, 16) -- 12829
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(12,12)), 0, 16) -- 12830
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(13,13)), 0, 16) -- 12831
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(14,14)), 0, 16) -- 12832
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(15,15)), 0, 16) -- 12833
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(16,16)), 0, 16) -- 12834
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(17,17)), 0, 16) -- 12835
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),( 9, 9)), 0, 16) -- 12836
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(10,10)), 0, 16) -- 12837
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(11,11)), 0, 16) -- 12838
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(12,12)), 0, 16) -- 12839
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(13,13)), 0, 16) -- 12840
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(14,14)), 0, 16) -- 12841
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(15,15)), 0, 16) -- 12842
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(16,16)), 0, 16) -- 12843
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 12844
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 12845
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 12846
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 12847
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 12848
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 12849
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 12850
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 12851
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 12852
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 12853
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 12854
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 12855
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 12856
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 12857
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 12858
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 12859
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(19,19),(11,11)), 0, 15) -- 12860
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(20,20),(12,12)), 0, 15) -- 12861
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(21,21),(13,13)), 0, 15) -- 12862
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(22,22),(14,14)), 0, 15) -- 12863
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(23,23),(15,15)), 0, 15) -- 12864
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(24,24),(16,16)), 0, 15) -- 12865
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(25,25),(17,17)), 0, 15) -- 12866
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(26,26),(18,18)), 0, 15) -- 12867
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(19,19),(12,12)), 0, 15) -- 12868
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(20,20),(13,13)), 0, 15) -- 12869
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(21,21),(14,14)), 0, 15) -- 12870
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(22,22),(15,15)), 0, 15) -- 12871
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(23,23),(16,16)), 0, 15) -- 12872
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(24,24),(17,17)), 0, 15) -- 12873
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(25,25),(18,18)), 0, 15) -- 12874
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(26,26),(19,19)), 0, 15) -- 12875
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(19,19),(10,10)), 0, 15) -- 12876
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(20,20),(11,11)), 0, 15) -- 12877
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(21,21),(12,12)), 0, 15) -- 12878
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(22,22),(13,13)), 0, 15) -- 12879
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(23,23),(14,14)), 0, 15) -- 12880
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(24,24),(15,15)), 0, 15) -- 12881
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(25,25),(16,16)), 0, 15) -- 12882
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(26,26),(17,17)), 0, 15) -- 12883
,( 10, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(10,10)), 0, 15) -- 12884
,( 10, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(11,11)), 0, 15) -- 12885
,( 10, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(12,12)), 0, 15) -- 12886
,( 10, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(13,13)), 0, 15) -- 12887
,( 10, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(14,14)), 0, 15) -- 12888
,( 10, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(15,15)), 0, 15) -- 12889
,( 10, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(16,16)), 0, 15) -- 12890
,( 10, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(17,17)), 0, 15) -- 12891
,( 10, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 12892
,( 10, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 12893
,( 10, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 12894
,( 10, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 12895
,( 10, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 12896
,( 10, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 12897
,( 10, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 12898
,( 10, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 12899
,( 10, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 12900
,( 10, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 12901
,( 10, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 12902
,( 10, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 12903
,( 10, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 12904
,( 10, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 12905
,( 10, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 12906
,( 10, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 12907
,( 10, E,0,0,((26,29),(22,23),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 12908
,( 10, E,0,0,((28,31),(24,25),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 12909
,( 10, E,0,0,((30,33),(26,27),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 12910
,( 10, E,0,0,((32,35),(28,29),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 12911
,( 10, E,0,0,((26,29),(22,23),( 0, 1),(17,17),(20,20),(10,13)), 0, 14) -- 12912
,( 10, E,0,0,((28,31),(24,25),( 2, 3),(19,19),(22,22),(12,15)), 0, 14) -- 12913
,( 10, E,0,0,((30,33),(26,27),( 4, 5),(21,21),(24,24),(14,17)), 0, 14) -- 12914
,( 10, E,0,0,((32,35),(28,29),( 6, 7),(23,23),(26,26),(16,19)), 0, 14) -- 12915
,( 10, E,0,0,((26,29),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 14) -- 12916
,( 10, E,0,0,((28,31),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 14) -- 12917
,( 10, E,0,0,((30,33),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 14) -- 12918
,( 10, E,0,0,((32,35),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 14) -- 12919
,( 10, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),( 8,11)), 0, 14) -- 12920
,( 10, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(10,13)), 0, 14) -- 12921
,( 10, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(12,15)), 0, 14) -- 12922
,( 10, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(14,17)), 0, 14) -- 12923
,( 10, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(12,15)), 0, 13) -- 12924
,( 10, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(14,17)), 0, 13) -- 12925
,( 10, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(16,19)), 0, 13) -- 12926
,( 10, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(18,21)), 0, 13) -- 12927
,( 10, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(10,13)), 0, 13) -- 12928
,( 10, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(12,15)), 0, 13) -- 12929
,( 10, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(14,17)), 0, 13) -- 12930
,( 10, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(16,19)), 0, 13) -- 12931
,( 10, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 12932
,( 10, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 12933
,( 10, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 12934
,( 10, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 12935
,( 10, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,20),( 8,11)), 0, 12) -- 12936
,( 10, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,22),(10,13)), 0, 12) -- 12937
,( 10, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,24),(12,15)), 0, 12) -- 12938
,( 10, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,26),(14,17)), 0, 12) -- 12939
,( 10, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 12) -- 12940
,( 10, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 12) -- 12941
,( 10, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 12) -- 12942
,( 10, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 12) -- 12943
,( 10, E,0,0,((26,29),(22,22),( 1, 1),(18,19),(22,22),(14,17)), 0, 12) -- 12944
,( 10, E,0,0,((28,31),(24,24),( 3, 3),(20,21),(24,24),(16,19)), 0, 12) -- 12945
,( 10, E,0,0,((30,33),(26,26),( 5, 5),(22,23),(26,26),(18,21)), 0, 12) -- 12946
,( 10, E,0,0,((32,35),(28,28),( 7, 7),(24,25),(28,28),(20,23)), 0, 12) -- 12947
,( 10, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 11) -- 12948
,( 10, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 11) -- 12949
,( 10, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 11) -- 12950
,( 10, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 11) -- 12951
,( 10, E,0,0,((24,27),(20,21),( 0, 0),(16,17),(18,19),( 8,11)), 0, 11) -- 12952
,( 10, E,0,0,((26,29),(22,23),( 2, 2),(18,19),(20,21),(10,13)), 0, 11) -- 12953
,( 10, E,0,0,((28,31),(24,25),( 4, 4),(20,21),(22,23),(12,15)), 0, 11) -- 12954
,( 10, E,0,0,((30,33),(26,27),( 6, 6),(22,23),(24,25),(14,17)), 0, 11) -- 12955
,( 10, E,0,0,((24,27),(20,21),( 1, 1),(18,19),(22,23),(10,13)), 0, 11) -- 12956
,( 10, E,0,0,((26,29),(22,23),( 3, 3),(20,21),(24,25),(12,15)), 0, 11) -- 12957
,( 10, E,0,0,((28,31),(24,25),( 5, 5),(22,23),(26,27),(14,17)), 0, 11) -- 12958
,( 10, E,0,0,((30,33),(26,27),( 7, 7),(24,25),(28,29),(16,19)), 0, 11) -- 12959
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 12960
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 12961
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 12962
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 12963
,( 10, E,0,0,((22,25),(19,19),( 0, 0),(18,19),(20,21),(10,13)), 0, 10) -- 12964
,( 10, E,0,0,((24,27),(21,21),( 2, 2),(20,21),(22,23),(12,15)), 0, 10) -- 12965
,( 10, E,0,0,((26,29),(23,23),( 4, 4),(22,23),(24,25),(14,17)), 0, 10) -- 12966
,( 10, E,0,0,((28,31),(25,25),( 6, 6),(24,25),(26,27),(16,19)), 0, 10) -- 12967
,( 10, E,0,0,((22,25),(20,20),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 12968
,( 10, E,0,0,((24,27),(22,22),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 12969
,( 10, E,0,0,((26,29),(24,24),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 12970
,( 10, E,0,0,((28,31),(26,26),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 12971
,( 10, E,0,0,((22,25),(19,19),( 0, 0),(17,17),(20,21),(10,13)), 0, 10) -- 12972
,( 10, E,0,0,((24,27),(21,21),( 2, 2),(19,19),(22,23),(12,15)), 0, 10) -- 12973
,( 10, E,0,0,((26,29),(23,23),( 4, 4),(21,21),(24,25),(14,17)), 0, 10) -- 12974
,( 10, E,0,0,((28,31),(25,25),( 6, 6),(23,23),(26,27),(16,19)), 0, 10) -- 12975
,( 10, E,0,0,((23,23),(20,20),( 0, 1),(18,19),(20,21),(10,13)), 0, 10) -- 12976
,( 10, E,0,0,((25,25),(22,22),( 2, 3),(20,21),(22,23),(12,15)), 0, 10) -- 12977
,( 10, E,0,0,((27,27),(24,24),( 4, 5),(22,23),(24,25),(14,17)), 0, 10) -- 12978
,( 10, E,0,0,((29,29),(26,26),( 6, 7),(24,25),(26,27),(16,19)), 0, 10) -- 12979
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(16,19)), 0, 10) -- 12980
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(18,21)), 0, 10) -- 12981
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(20,23)), 0, 10) -- 12982
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(22,23)), 0, 10) -- 12983
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0, 10) -- 12984
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0, 10) -- 12985
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0, 10) -- 12986
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0, 10) -- 12987
,( 10, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(24,24),(14,17)), 0, 10) -- 12988
,( 10, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(26,26),(16,19)), 0, 10) -- 12989
,( 10, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(28,28),(18,21)), 0, 10) -- 12990
,( 10, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(30,30),(20,23)), 0, 10) -- 12991
,( 10, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(12,15)), 0, 10) -- 12992
,( 10, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(14,17)), 0, 10) -- 12993
,( 10, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(16,19)), 0, 10) -- 12994
,( 10, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(18,21)), 0, 10) -- 12995
,( 10, E,0,0,((22,25),(20,21),( 1, 1),(19,19),(24,24),(16,19)), 0, 10) -- 12996
,( 10, E,0,0,((24,27),(22,23),( 3, 3),(21,21),(26,26),(18,21)), 0, 10) -- 12997
,( 10, E,0,0,((26,29),(24,25),( 5, 5),(23,23),(28,28),(20,23)), 0, 10) -- 12998
,( 10, E,0,0,((28,31),(26,27),( 7, 7),(25,25),(30,30),(22,23)), 0, 10) -- 12999
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 8,11)), 0,  9) -- 13000
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(10,13)), 0,  9) -- 13001
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(12,15)), 0,  9) -- 13002
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(14,17)), 0,  9) -- 13003
,( 10, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 13004
,( 10, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 13005
,( 10, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 13006
,( 10, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 13007
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(20,21),(24,25),(12,15)), 0,  9) -- 13008
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(22,23),(26,27),(14,17)), 0,  9) -- 13009
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(24,25),(28,29),(16,19)), 0,  9) -- 13010
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(26,27),(30,31),(18,21)), 0,  9) -- 13011
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(18,19),( 4, 5)), 0,  9) -- 13012
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(20,21),( 6, 7)), 0,  9) -- 13013
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(22,23),( 8, 9)), 0,  9) -- 13014
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(24,25),(10,11)), 0,  9) -- 13015
,( 10, E,0,0,((22,25),(20,20),( 1, 1),(18,19),(22,23),( 8,11)), 0,  9) -- 13016
,( 10, E,0,0,((24,27),(22,22),( 3, 3),(20,21),(24,25),(10,13)), 0,  9) -- 13017
,( 10, E,0,0,((26,29),(24,24),( 5, 5),(22,23),(26,27),(12,15)), 0,  9) -- 13018
,( 10, E,0,0,((28,31),(26,26),( 7, 7),(24,25),(28,29),(14,17)), 0,  9) -- 13019
,( 10, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 13020
,( 10, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 13021
,( 10, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 13022
,( 10, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 13023
,( 10, E,0,0,((18,21),(18,19),( 0, 0),(18,19),(21,21),(10,13)), 0,  9) -- 13024
,( 10, E,0,0,((20,23),(20,21),( 2, 2),(20,21),(23,23),(12,15)), 0,  9) -- 13025
,( 10, E,0,0,((22,25),(22,23),( 4, 4),(22,23),(25,25),(14,17)), 0,  9) -- 13026
,( 10, E,0,0,((24,27),(24,25),( 6, 6),(24,25),(27,27),(16,19)), 0,  9) -- 13027
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 2, 5)), 0,  9) -- 13028
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 4, 7)), 0,  9) -- 13029
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),( 6, 9)), 0,  9) -- 13030
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),( 8,11)), 0,  9) -- 13031
,( 10, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 13032
,( 10, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 13033
,( 10, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 13034
,( 10, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 13035
,( 10, E,0,0,((18,21),(17,17),( 0, 0),(18,19),(22,23),(10,13)), 0,  9) -- 13036
,( 10, E,0,0,((20,23),(19,19),( 2, 2),(20,21),(24,25),(12,15)), 0,  9) -- 13037
,( 10, E,0,0,((22,25),(21,21),( 4, 4),(22,23),(26,27),(14,17)), 0,  9) -- 13038
,( 10, E,0,0,((24,27),(23,23),( 6, 6),(24,25),(28,29),(16,19)), 0,  9) -- 13039
,( 10, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(19,19),( 4, 7)), 0,  9) -- 13040
,( 10, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(21,21),( 6, 9)), 0,  9) -- 13041
,( 10, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(23,23),( 8,11)), 0,  9) -- 13042
,( 10, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(25,25),(10,13)), 0,  9) -- 13043
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(19,19),(24,25),(14,17)), 0,  9) -- 13044
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(21,21),(26,27),(16,19)), 0,  9) -- 13045
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(23,23),(28,29),(18,21)), 0,  9) -- 13046
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(25,25),(30,31),(20,23)), 0,  9) -- 13047
,( 10, E,0,0,((20,23),(18,19),( 0, 0),(17,17),(18,19),( 4, 7)), 0,  9) -- 13048
,( 10, E,0,0,((22,25),(20,21),( 2, 2),(19,19),(20,21),( 6, 9)), 0,  9) -- 13049
,( 10, E,0,0,((24,27),(22,23),( 4, 4),(21,21),(22,23),( 8,11)), 0,  9) -- 13050
,( 10, E,0,0,((26,29),(24,25),( 6, 6),(23,23),(24,25),(10,13)), 0,  9) -- 13051
,( 10, E,0,0,((20,23),(18,19),( 0, 1),(20,20),(24,25),(16,19)), 0,  9) -- 13052
,( 10, E,0,0,((22,25),(20,21),( 2, 3),(22,22),(26,27),(18,21)), 0,  9) -- 13053
,( 10, E,0,0,((24,27),(22,23),( 4, 5),(24,24),(28,29),(20,23)), 0,  9) -- 13054
,( 10, E,0,0,((26,29),(24,25),( 6, 7),(26,26),(30,31),(22,23)), 0,  9) -- 13055
,( 10, E,0,0,((16,19),(16,17),( 0, 0),(19,19),(24,25),(12,15)), 0,  9) -- 13056
,( 10, E,0,0,((18,21),(18,19),( 2, 2),(21,21),(26,27),(14,17)), 0,  9) -- 13057
,( 10, E,0,0,((20,23),(20,21),( 4, 4),(23,23),(28,29),(16,19)), 0,  9) -- 13058
,( 10, E,0,0,((22,25),(22,23),( 6, 6),(25,25),(30,31),(18,21)), 0,  9) -- 13059
,( 10, E,0,0,((18,21),(18,19),( 0, 0),(18,19),(22,23),( 6, 9)), 0,  9) -- 13060
,( 10, E,0,0,((20,23),(20,21),( 2, 2),(20,21),(24,25),( 8,11)), 0,  9) -- 13061
,( 10, E,0,0,((22,25),(22,23),( 4, 4),(22,23),(26,27),(10,13)), 0,  9) -- 13062
,( 10, E,0,0,((24,27),(24,25),( 6, 6),(24,25),(28,29),(12,15)), 0,  9) -- 13063
,( 10, E,0,0,((18,21),(18,19),( 1, 1),(20,21),(26,27),(16,19)), 0,  9) -- 13064
,( 10, E,0,0,((20,23),(20,21),( 3, 3),(22,23),(28,29),(18,21)), 0,  9) -- 13065
,( 10, E,0,0,((22,25),(22,23),( 5, 5),(24,25),(30,31),(20,23)), 0,  9) -- 13066
,( 10, E,0,0,((24,27),(24,25),( 7, 7),(26,27),(32,33),(22,23)), 0,  9) -- 13067
,( 10, E,0,0,((20,23),(19,19),( 1, 1),(20,20),(22,23),(12,15)), 0,  9) -- 13068
,( 10, E,0,0,((22,25),(21,21),( 3, 3),(22,22),(24,25),(14,17)), 0,  9) -- 13069
,( 10, E,0,0,((24,27),(23,23),( 5, 5),(24,24),(26,27),(16,19)), 0,  9) -- 13070
,( 10, E,0,0,((26,29),(25,25),( 7, 7),(26,26),(28,29),(18,21)), 0,  9) -- 13071
,( 10, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(22,25),( 8,11)), 0,  8) -- 13072
,( 10, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(24,27),(10,13)), 0,  8) -- 13073
,( 10, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(26,29),(12,15)), 0,  8) -- 13074
,( 10, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(28,31),(14,17)), 0,  8) -- 13075
,( 10, E,0,0,((18,21),(16,19),( 0, 1),(18,21),(18,21),( 0, 0)), 0,  8) -- 13076
,( 10, E,0,0,((20,23),(18,21),( 2, 3),(20,23),(20,23),( 2, 2)), 0,  8) -- 13077
,( 10, E,0,0,((22,25),(20,23),( 4, 5),(22,25),(22,25),( 4, 4)), 0,  8) -- 13078
,( 10, E,0,0,((24,27),(22,25),( 6, 7),(24,27),(24,27),( 6, 6)), 0,  8) -- 13079
,( 10, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(16,19),( 2, 3)), 0,  8) -- 13080
,( 10, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(18,21),( 4, 5)), 0,  8) -- 13081
,( 10, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(20,23),( 6, 7)), 0,  8) -- 13082
,( 10, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(22,25),( 8, 9)), 0,  8) -- 13083
,( 10, E,0,0,((14,17),(14,17),( 0, 1),(18,21),(18,21),(99,99)), 0,  7) -- 13084
,( 10, E,0,0,((16,19),(16,19),( 2, 3),(20,23),(20,23),(99,99)), 0,  7) -- 13085
,( 10, E,0,0,((18,21),(18,21),( 4, 5),(22,25),(22,25),(99,99)), 0,  7) -- 13086
,( 10, E,0,0,((20,23),(20,23),( 6, 7),(24,27),(24,27),(99,99)), 0,  7) -- 13087
,( 10, E,0,0,((16,19),(16,19),( 0, 1),(16,19),(14,17),(99,99)), 0,  7) -- 13088
,( 10, E,0,0,((18,21),(18,21),( 2, 3),(18,21),(16,19),(99,99)), 0,  7) -- 13089
,( 10, E,0,0,((20,23),(20,23),( 4, 5),(20,23),(18,21),(99,99)), 0,  7) -- 13090
,( 10, E,0,0,((22,25),(22,25),( 6, 7),(22,25),(20,23),(99,99)), 0,  7) -- 13091
,( 10, E,0,0,((14,17),(14,17),( 0, 1),(18,21),(22,25),(99,99)), 0,  7) -- 13092
,( 10, E,0,0,((16,19),(16,19),( 2, 3),(20,23),(24,27),(99,99)), 0,  7) -- 13093
,( 10, E,0,0,((18,21),(18,21),( 4, 5),(22,25),(26,29),(99,99)), 0,  7) -- 13094
,( 10, E,0,0,((20,23),(20,23),( 6, 7),(24,27),(28,31),(99,99)), 0,  7) -- 13095
,( 10, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 13096
,( 10, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 13097
,( 10, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 13098
,( 10, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 13099
,( 10, E,0,1,((16,19),(16,19),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 13100
,( 10, E,0,1,((18,21),(18,21),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 13101
,( 10, E,0,1,((20,23),(20,23),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 13102
,( 10, E,0,1,((22,25),(22,25),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 13103
,( 10, E,0,1,(( 8,11),(12,15),( 0, 1),(18,21),(99,99),(99,99)), 0,  6) -- 13104
,( 10, E,0,1,((10,13),(14,17),( 2, 3),(20,23),(99,99),(99,99)), 0,  6) -- 13105
,( 10, E,0,1,((12,15),(16,19),( 4, 5),(22,25),(99,99),(99,99)), 0,  6) -- 13106
,( 10, E,0,1,((14,17),(18,21),( 6, 7),(24,27),(99,99),(99,99)), 0,  6) -- 13107
,( 10, E,0,1,((12,15),(14,17),( 0, 1),(14,17),(99,99),(99,99)), 0,  6) -- 13108
,( 10, E,0,1,((14,17),(16,19),( 2, 3),(16,19),(99,99),(99,99)), 0,  6) -- 13109
,( 10, E,0,1,((16,19),(18,21),( 4, 5),(18,21),(99,99),(99,99)), 0,  6) -- 13110
,( 10, E,0,1,((18,21),(20,23),( 6, 7),(20,23),(99,99),(99,99)), 0,  6) -- 13111
,( 10, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 13112
,( 10, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 13113
,( 10, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 13114
,( 10, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 13115
,( 10, E,0,1,(( 4, 7),(12,15),( 0, 1),(16,19),(99,99),(99,99)), 0,  5) -- 13116
,( 10, E,0,1,(( 6, 9),(14,17),( 2, 3),(18,21),(99,99),(99,99)), 0,  5) -- 13117
,( 10, E,0,1,(( 8,11),(16,19),( 4, 5),(20,23),(99,99),(99,99)), 0,  5) -- 13118
,( 10, E,0,1,((10,13),(18,21),( 6, 7),(22,25),(99,99),(99,99)), 0,  5) -- 13119
,( 10, E,0,1,((20,23),(20,23),( 0, 1),(10,13),(99,99),(99,99)), 0,  5) -- 13120
,( 10, E,0,1,((22,25),(22,25),( 2, 3),(12,15),(99,99),(99,99)), 0,  5) -- 13121
,( 10, E,0,1,((24,27),(24,27),( 4, 5),(14,17),(99,99),(99,99)), 0,  5) -- 13122
,( 10, E,0,1,((26,29),(26,29),( 6, 7),(16,19),(99,99),(99,99)), 0,  5) -- 13123
,( 10, E,0,1,(( 4, 5),(10,13),( 0, 1),(18,21),(99,99),(99,99)), 0,  5) -- 13124
,( 10, E,0,1,(( 6, 7),(12,15),( 2, 3),(20,23),(99,99),(99,99)), 0,  5) -- 13125
,( 10, E,0,1,(( 8, 9),(14,17),( 4, 5),(22,25),(99,99),(99,99)), 0,  5) -- 13126
,( 10, E,0,1,((10,11),(16,19),( 6, 7),(24,27),(99,99),(99,99)), 0,  5) -- 13127
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 13128
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 13129
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 13130
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 13131
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 13132
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 13133
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 13134
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 13135
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 13136
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 13137
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 13138
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 13139
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 13140
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 13141
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 13142
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 13143
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(16,16),( 7, 7)), 1, 31) -- 13144
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(17,17),( 8, 8)), 1, 31) -- 13145
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(18,18),( 9, 9)), 1, 31) -- 13146
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(19,19),(10,10)), 1, 31) -- 13147
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(20,20),(11,11)), 1, 31) -- 13148
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(21,21),(12,12)), 1, 31) -- 13149
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(22,22),(13,13)), 1, 31) -- 13150
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(23,23),(14,14)), 1, 31) -- 13151
,( 11, E,0,0,((32,32),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 31) -- 13152
,( 11, E,0,0,((33,33),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 31) -- 13153
,( 11, E,0,0,((34,34),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 31) -- 13154
,( 11, E,0,0,((35,35),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 31) -- 13155
,( 11, E,0,0,((36,36),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 31) -- 13156
,( 11, E,0,0,((37,37),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 31) -- 13157
,( 11, E,0,0,((38,38),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 31) -- 13158
,( 11, E,0,0,((39,39),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 31) -- 13159
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 31) -- 13160
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 31) -- 13161
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 31) -- 13162
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 31) -- 13163
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 31) -- 13164
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 31) -- 13165
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 31) -- 13166
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 31) -- 13167
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 1, 31) -- 13168
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 1, 31) -- 13169
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 1, 31) -- 13170
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 1, 31) -- 13171
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 1, 31) -- 13172
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 1, 31) -- 13173
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 1, 31) -- 13174
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 1, 31) -- 13175
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 8, 8)), 1, 31) -- 13176
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 9, 9)), 1, 31) -- 13177
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),(10,10)), 1, 31) -- 13178
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),(11,11)), 1, 31) -- 13179
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(12,12)), 1, 31) -- 13180
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(13,13)), 1, 31) -- 13181
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(14,14)), 1, 31) -- 13182
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(15,15)), 1, 31) -- 13183
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 30) -- 13184
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 30) -- 13185
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),(10,10)), 1, 30) -- 13186
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(11,11)), 1, 30) -- 13187
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(12,12)), 1, 30) -- 13188
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(13,13)), 1, 30) -- 13189
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(14,14)), 1, 30) -- 13190
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(15,15)), 1, 30) -- 13191
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(16,16),( 7, 7)), 1, 26) -- 13192
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(17,17),( 8, 8)), 1, 26) -- 13193
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(18,18),( 9, 9)), 1, 26) -- 13194
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(19,19),(10,10)), 1, 26) -- 13195
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(20,20),(11,11)), 1, 26) -- 13196
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(21,21),(12,12)), 1, 26) -- 13197
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(22,22),(13,13)), 1, 26) -- 13198
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(23,23),(14,14)), 1, 26) -- 13199
,( 11, E,0,0,((33,33),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 1, 25) -- 13200
,( 11, E,0,0,((34,34),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 1, 25) -- 13201
,( 11, E,0,0,((35,35),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 1, 25) -- 13202
,( 11, E,0,0,((36,36),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 1, 25) -- 13203
,( 11, E,0,0,((37,37),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 1, 25) -- 13204
,( 11, E,0,0,((38,38),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 1, 25) -- 13205
,( 11, E,0,0,((39,39),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 1, 25) -- 13206
,( 11, E,0,0,((40,40),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 1, 25) -- 13207
,( 11, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 13208
,( 11, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 13209
,( 11, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 13210
,( 11, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 13211
,( 11, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 13212
,( 11, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 13213
,( 11, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 13214
,( 11, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 13215
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 24) -- 13216
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 24) -- 13217
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 24) -- 13218
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 24) -- 13219
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 24) -- 13220
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 24) -- 13221
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 24) -- 13222
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 24) -- 13223
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 23) -- 13224
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 23) -- 13225
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 23) -- 13226
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 23) -- 13227
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 23) -- 13228
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 23) -- 13229
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 23) -- 13230
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 23) -- 13231
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 23) -- 13232
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 23) -- 13233
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 23) -- 13234
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 23) -- 13235
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 23) -- 13236
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 23) -- 13237
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 23) -- 13238
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 23) -- 13239
,( 11, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 21) -- 13240
,( 11, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 21) -- 13241
,( 11, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 21) -- 13242
,( 11, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 21) -- 13243
,( 11, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(19,19),(10,10)), 1, 21) -- 13244
,( 11, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(20,20),(11,11)), 1, 21) -- 13245
,( 11, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(21,21),(12,12)), 1, 21) -- 13246
,( 11, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(22,22),(13,13)), 1, 21) -- 13247
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 20) -- 13248
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 20) -- 13249
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 20) -- 13250
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 20) -- 13251
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 20) -- 13252
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 20) -- 13253
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 20) -- 13254
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 20) -- 13255
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(16,16),(15,15),( 7, 7)), 1, 20) -- 13256
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(17,17),(16,16),( 8, 8)), 1, 20) -- 13257
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(18,18),(17,17),( 9, 9)), 1, 20) -- 13258
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(19,19),(18,18),(10,10)), 1, 20) -- 13259
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(20,20),(19,19),(11,11)), 1, 20) -- 13260
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(21,21),(20,20),(12,12)), 1, 20) -- 13261
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(22,22),(21,21),(13,13)), 1, 20) -- 13262
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(23,23),(22,22),(14,14)), 1, 20) -- 13263
,( 11, E,0,0,((33,33),(24,24),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 20) -- 13264
,( 11, E,0,0,((34,34),(25,25),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 20) -- 13265
,( 11, E,0,0,((35,35),(26,26),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 20) -- 13266
,( 11, E,0,0,((36,36),(27,27),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 20) -- 13267
,( 11, E,0,0,((37,37),(28,28),( 4, 4),(19,19),(18,18),(10,10)), 1, 20) -- 13268
,( 11, E,0,0,((38,38),(29,29),( 5, 5),(20,20),(19,19),(11,11)), 1, 20) -- 13269
,( 11, E,0,0,((39,39),(30,30),( 6, 6),(21,21),(20,20),(12,12)), 1, 20) -- 13270
,( 11, E,0,0,((40,40),(31,31),( 7, 7),(22,22),(21,21),(13,13)), 1, 20) -- 13271
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 20) -- 13272
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 20) -- 13273
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 20) -- 13274
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),(10,10)), 1, 20) -- 13275
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(11,11)), 1, 20) -- 13276
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(12,12)), 1, 20) -- 13277
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(13,13)), 1, 20) -- 13278
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(14,14)), 1, 20) -- 13279
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 19) -- 13280
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 19) -- 13281
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 19) -- 13282
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 19) -- 13283
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(19,19),(10,10)), 1, 19) -- 13284
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(20,20),(11,11)), 1, 19) -- 13285
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(21,21),(12,12)), 1, 19) -- 13286
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(22,22),(13,13)), 1, 19) -- 13287
,( 11, E,0,0,((33,33),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 19) -- 13288
,( 11, E,0,0,((34,34),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 19) -- 13289
,( 11, E,0,0,((35,35),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 19) -- 13290
,( 11, E,0,0,((36,36),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 19) -- 13291
,( 11, E,0,0,((37,37),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 19) -- 13292
,( 11, E,0,0,((38,38),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 19) -- 13293
,( 11, E,0,0,((39,39),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 19) -- 13294
,( 11, E,0,0,((40,40),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 19) -- 13295
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 18) -- 13296
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 18) -- 13297
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 18) -- 13298
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 18) -- 13299
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 18) -- 13300
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 18) -- 13301
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 18) -- 13302
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 18) -- 13303
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 18) -- 13304
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 18) -- 13305
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 18) -- 13306
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 18) -- 13307
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 18) -- 13308
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 18) -- 13309
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 18) -- 13310
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 18) -- 13311
,( 11, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 18) -- 13312
,( 11, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 18) -- 13313
,( 11, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 18) -- 13314
,( 11, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 18) -- 13315
,( 11, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 18) -- 13316
,( 11, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 18) -- 13317
,( 11, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 18) -- 13318
,( 11, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 18) -- 13319
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 18) -- 13320
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 18) -- 13321
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 18) -- 13322
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 18) -- 13323
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 18) -- 13324
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 18) -- 13325
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 18) -- 13326
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 18) -- 13327
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 6, 6)), 1, 17) -- 13328
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 7, 7)), 1, 17) -- 13329
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 8, 8)), 1, 17) -- 13330
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),( 9, 9)), 1, 17) -- 13331
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(10,10)), 1, 17) -- 13332
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(11,11)), 1, 17) -- 13333
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(12,12)), 1, 17) -- 13334
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(13,13)), 1, 17) -- 13335
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 17) -- 13336
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 17) -- 13337
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 17) -- 13338
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 17) -- 13339
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),(10,10)), 1, 17) -- 13340
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(11,11)), 1, 17) -- 13341
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(12,12)), 1, 17) -- 13342
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(13,13)), 1, 17) -- 13343
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 17) -- 13344
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 17) -- 13345
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 17) -- 13346
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 17) -- 13347
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 17) -- 13348
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 17) -- 13349
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 17) -- 13350
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 17) -- 13351
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 17) -- 13352
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 17) -- 13353
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 17) -- 13354
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 17) -- 13355
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 17) -- 13356
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 17) -- 13357
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 17) -- 13358
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 17) -- 13359
,( 11, E,0,0,((34,34),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 17) -- 13360
,( 11, E,0,0,((35,35),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 17) -- 13361
,( 11, E,0,0,((36,36),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 17) -- 13362
,( 11, E,0,0,((37,37),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 17) -- 13363
,( 11, E,0,0,((38,38),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 17) -- 13364
,( 11, E,0,0,((39,39),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 17) -- 13365
,( 11, E,0,0,((40,40),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 17) -- 13366
,( 11, E,0,0,((41,41),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 17) -- 13367
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(15,15),(15,15),( 7, 7)), 1, 16) -- 13368
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(16,16),(16,16),( 8, 8)), 1, 16) -- 13369
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(17,17),(17,17),( 9, 9)), 1, 16) -- 13370
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(18,18),(18,18),(10,10)), 1, 16) -- 13371
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(19,19),(19,19),(11,11)), 1, 16) -- 13372
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(20,20),(20,20),(12,12)), 1, 16) -- 13373
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(21,21),(21,21),(13,13)), 1, 16) -- 13374
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(22,22),(22,22),(14,14)), 1, 16) -- 13375
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 16) -- 13376
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 16) -- 13377
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 16) -- 13378
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 16) -- 13379
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 16) -- 13380
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(10,10)), 1, 16) -- 13381
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(11,11)), 1, 16) -- 13382
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(12,12)), 1, 16) -- 13383
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(15,15),(14,14),( 6, 6)), 1, 16) -- 13384
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(16,16),(15,15),( 7, 7)), 1, 16) -- 13385
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(17,17),(16,16),( 8, 8)), 1, 16) -- 13386
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(18,18),(17,17),( 9, 9)), 1, 16) -- 13387
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(19,19),(18,18),(10,10)), 1, 16) -- 13388
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(20,20),(19,19),(11,11)), 1, 16) -- 13389
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(21,21),(20,20),(12,12)), 1, 16) -- 13390
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(22,22),(21,21),(13,13)), 1, 16) -- 13391
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 13392
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 13393
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 13394
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 13395
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 13396
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 13397
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 13398
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 13399
,( 11, E,0,0,((36,36),(26,26),( 0, 0),(15,15),(14,14),( 5, 5)), 1, 15) -- 13400
,( 11, E,0,0,((37,37),(27,27),( 1, 1),(16,16),(15,15),( 6, 6)), 1, 15) -- 13401
,( 11, E,0,0,((38,38),(28,28),( 2, 2),(17,17),(16,16),( 7, 7)), 1, 15) -- 13402
,( 11, E,0,0,((39,39),(29,29),( 3, 3),(18,18),(17,17),( 8, 8)), 1, 15) -- 13403
,( 11, E,0,0,((40,40),(30,30),( 4, 4),(19,19),(18,18),( 9, 9)), 1, 15) -- 13404
,( 11, E,0,0,((41,41),(31,31),( 5, 5),(20,20),(19,19),(10,10)), 1, 15) -- 13405
,( 11, E,0,0,((42,42),(32,32),( 6, 6),(21,21),(20,20),(11,11)), 1, 15) -- 13406
,( 11, E,0,0,((43,43),(33,33),( 7, 7),(22,22),(21,21),(12,12)), 1, 15) -- 13407
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 13408
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 13409
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 13410
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 13411
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 13412
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 13413
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 13414
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 13415
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(13,13),( 4, 4)), 1, 15) -- 13416
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(14,14),( 5, 5)), 1, 15) -- 13417
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(15,15),( 6, 6)), 1, 15) -- 13418
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(16,16),( 7, 7)), 1, 15) -- 13419
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(17,17),( 8, 8)), 1, 15) -- 13420
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(18,18),( 9, 9)), 1, 15) -- 13421
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(19,19),(10,10)), 1, 15) -- 13422
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(20,20),(11,11)), 1, 15) -- 13423
,( 11, E,0,0,((35,35),(26,26),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 13424
,( 11, E,0,0,((36,36),(27,27),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 13425
,( 11, E,0,0,((37,37),(28,28),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 13426
,( 11, E,0,0,((38,38),(29,29),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 13427
,( 11, E,0,0,((39,39),(30,30),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 13428
,( 11, E,0,0,((40,40),(31,31),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 13429
,( 11, E,0,0,((41,41),(32,32),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 13430
,( 11, E,0,0,((42,42),(33,33),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 13431
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 6, 6)), 1, 15) -- 13432
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 7, 7)), 1, 15) -- 13433
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 8, 8)), 1, 15) -- 13434
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 9, 9)), 1, 15) -- 13435
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),(10,10)), 1, 15) -- 13436
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(11,11)), 1, 15) -- 13437
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(12,12)), 1, 15) -- 13438
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(13,13)), 1, 15) -- 13439
,( 11, E,0,0,((34,34),(25,25),( 0, 0),(14,14),(13,13),( 5, 5)), 1, 15) -- 13440
,( 11, E,0,0,((35,35),(26,26),( 1, 1),(15,15),(14,14),( 6, 6)), 1, 15) -- 13441
,( 11, E,0,0,((36,36),(27,27),( 2, 2),(16,16),(15,15),( 7, 7)), 1, 15) -- 13442
,( 11, E,0,0,((37,37),(28,28),( 3, 3),(17,17),(16,16),( 8, 8)), 1, 15) -- 13443
,( 11, E,0,0,((38,38),(29,29),( 4, 4),(18,18),(17,17),( 9, 9)), 1, 15) -- 13444
,( 11, E,0,0,((39,39),(30,30),( 5, 5),(19,19),(18,18),(10,10)), 1, 15) -- 13445
,( 11, E,0,0,((40,40),(31,31),( 6, 6),(20,20),(19,19),(11,11)), 1, 15) -- 13446
,( 11, E,0,0,((41,41),(32,32),( 7, 7),(21,21),(20,20),(12,12)), 1, 15) -- 13447
,( 11, E,0,0,((35,35),(25,25),( 0, 0),(14,14),(14,14),( 5, 5)), 1, 15) -- 13448
,( 11, E,0,0,((36,36),(26,26),( 1, 1),(15,15),(15,15),( 6, 6)), 1, 15) -- 13449
,( 11, E,0,0,((37,37),(27,27),( 2, 2),(16,16),(16,16),( 7, 7)), 1, 15) -- 13450
,( 11, E,0,0,((38,38),(28,28),( 3, 3),(17,17),(17,17),( 8, 8)), 1, 15) -- 13451
,( 11, E,0,0,((39,39),(29,29),( 4, 4),(18,18),(18,18),( 9, 9)), 1, 15) -- 13452
,( 11, E,0,0,((40,40),(30,30),( 5, 5),(19,19),(19,19),(10,10)), 1, 15) -- 13453
,( 11, E,0,0,((41,41),(31,31),( 6, 6),(20,20),(20,20),(11,11)), 1, 15) -- 13454
,( 11, E,0,0,((42,42),(32,32),( 7, 7),(21,21),(21,21),(12,12)), 1, 15) -- 13455
,( 11, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(14,15),( 4, 7)), 1, 14) -- 13456
,( 11, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(16,17),( 6, 9)), 1, 14) -- 13457
,( 11, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(18,19),( 8,11)), 1, 14) -- 13458
,( 11, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(20,21),(10,13)), 1, 14) -- 13459
,( 11, E,0,0,((34,37),(26,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 14) -- 13460
,( 11, E,0,0,((36,39),(28,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 14) -- 13461
,( 11, E,0,0,((38,41),(30,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 14) -- 13462
,( 11, E,0,0,((40,43),(32,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 14) -- 13463
,( 11, E,0,0,((36,39),(28,28),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 13) -- 13464
,( 11, E,0,0,((38,41),(30,30),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 13) -- 13465
,( 11, E,0,0,((40,43),(32,32),( 5, 5),(20,20),(18,19),( 8,11)), 1, 13) -- 13466
,( 11, E,0,0,((42,45),(34,34),( 7, 7),(22,22),(20,21),(10,13)), 1, 13) -- 13467
,( 11, E,0,0,((36,39),(27,27),( 1, 1),(16,16),(14,15),( 4, 7)), 1, 13) -- 13468
,( 11, E,0,0,((38,41),(29,29),( 3, 3),(18,18),(16,17),( 6, 9)), 1, 13) -- 13469
,( 11, E,0,0,((40,43),(31,31),( 5, 5),(20,20),(18,19),( 8,11)), 1, 13) -- 13470
,( 11, E,0,0,((42,45),(33,33),( 7, 7),(22,22),(20,21),(10,13)), 1, 13) -- 13471
,( 11, E,0,0,((36,39),(28,29),( 1, 1),(15,15),(14,14),( 4, 7)), 1, 13) -- 13472
,( 11, E,0,0,((38,41),(30,31),( 3, 3),(17,17),(16,16),( 6, 9)), 1, 13) -- 13473
,( 11, E,0,0,((40,43),(32,33),( 5, 5),(19,19),(18,18),( 8,11)), 1, 13) -- 13474
,( 11, E,0,0,((42,45),(34,35),( 7, 7),(21,21),(20,20),(10,13)), 1, 13) -- 13475
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 13476
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 13477
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 13478
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 13479
,( 11, E,0,0,((38,38),(27,27),( 0, 1),(14,15),(12,13),( 2, 5)), 1, 12) -- 13480
,( 11, E,0,0,((40,40),(29,29),( 2, 3),(16,17),(14,15),( 4, 7)), 1, 12) -- 13481
,( 11, E,0,0,((42,42),(31,31),( 4, 5),(18,19),(16,17),( 6, 9)), 1, 12) -- 13482
,( 11, E,0,0,((44,44),(33,33),( 6, 7),(20,21),(18,19),( 8,11)), 1, 12) -- 13483
,( 11, E,0,0,((36,39),(26,27),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 12) -- 13484
,( 11, E,0,0,((38,41),(28,29),( 2, 3),(16,17),(14,15),( 8,11)), 1, 12) -- 13485
,( 11, E,0,0,((40,43),(30,31),( 4, 5),(18,19),(16,17),(10,13)), 1, 12) -- 13486
,( 11, E,0,0,((42,45),(32,33),( 6, 7),(20,21),(18,19),(12,15)), 1, 12) -- 13487
,( 11, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(12,12),( 2, 5)), 1, 12) -- 13488
,( 11, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(14,14),( 4, 7)), 1, 12) -- 13489
,( 11, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(16,16),( 6, 9)), 1, 12) -- 13490
,( 11, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(18,18),( 8,11)), 1, 12) -- 13491
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(12,13),( 6, 9)), 1, 11) -- 13492
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(14,15),( 8,11)), 1, 11) -- 13493
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(16,17),(10,13)), 1, 11) -- 13494
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(18,19),(12,15)), 1, 11) -- 13495
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(12,13),(10,11),( 0, 3)), 1, 11) -- 13496
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(14,15),(12,13),( 2, 5)), 1, 11) -- 13497
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(16,17),(14,15),( 4, 7)), 1, 11) -- 13498
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(18,19),(16,17),( 6, 9)), 1, 11) -- 13499
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(11,11),( 0, 3)), 1, 11) -- 13500
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(13,13),( 2, 5)), 1, 11) -- 13501
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(15,15),( 4, 7)), 1, 11) -- 13502
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(17,17),( 6, 9)), 1, 11) -- 13503
,( 11, E,0,0,((36,39),(27,27),( 0, 0),(13,13),(10,11),( 0, 3)), 1, 11) -- 13504
,( 11, E,0,0,((38,41),(29,29),( 2, 2),(15,15),(12,13),( 2, 5)), 1, 11) -- 13505
,( 11, E,0,0,((40,43),(31,31),( 4, 4),(17,17),(14,15),( 4, 7)), 1, 11) -- 13506
,( 11, E,0,0,((42,45),(33,33),( 6, 6),(19,19),(16,17),( 6, 9)), 1, 11) -- 13507
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),( 6, 9)), 1, 11) -- 13508
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),( 8,11)), 1, 11) -- 13509
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(10,13)), 1, 11) -- 13510
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(12,15)), 1, 11) -- 13511
,( 11, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(12,13),( 2, 5)), 1, 10) -- 13512
,( 11, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(14,15),( 4, 7)), 1, 10) -- 13513
,( 11, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(16,17),( 6, 9)), 1, 10) -- 13514
,( 11, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(18,19),( 8,11)), 1, 10) -- 13515
,( 11, E,0,0,((38,41),(28,29),( 0, 0),(12,13),(12,13),( 4, 7)), 1, 10) -- 13516
,( 11, E,0,0,((40,43),(30,31),( 2, 2),(14,15),(14,15),( 6, 9)), 1, 10) -- 13517
,( 11, E,0,0,((42,45),(32,33),( 4, 4),(16,17),(16,17),( 8,11)), 1, 10) -- 13518
,( 11, E,0,0,((44,47),(34,35),( 6, 6),(18,19),(18,19),(10,13)), 1, 10) -- 13519
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(13,13),(10,11),( 4, 7)), 1, 10) -- 13520
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(15,15),(12,13),( 6, 9)), 1, 10) -- 13521
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(17,17),(14,15),( 8,11)), 1, 10) -- 13522
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(19,19),(16,17),(10,13)), 1, 10) -- 13523
,( 11, E,0,0,((42,45),(30,31),( 1, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 13524
,( 11, E,0,0,((44,47),(32,33),( 3, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 13525
,( 11, E,0,0,((46,49),(34,35),( 5, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 13526
,( 11, E,0,0,((48,51),(36,37),( 7, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 13527
,( 11, E,0,0,((40,43),(30,30),( 1, 1),(14,15),(12,13),( 6, 9)), 1, 10) -- 13528
,( 11, E,0,0,((42,45),(32,32),( 3, 3),(16,17),(14,15),( 8,11)), 1, 10) -- 13529
,( 11, E,0,0,((44,47),(34,34),( 5, 5),(18,19),(16,17),(10,13)), 1, 10) -- 13530
,( 11, E,0,0,((46,49),(36,36),( 7, 7),(20,21),(18,19),(12,15)), 1, 10) -- 13531
,( 11, E,0,0,((40,43),(29,29),( 0, 1),(14,14),(10,11),( 2, 5)), 1, 10) -- 13532
,( 11, E,0,0,((42,45),(31,31),( 2, 3),(16,16),(12,13),( 4, 7)), 1, 10) -- 13533
,( 11, E,0,0,((44,47),(33,33),( 4, 5),(18,18),(14,15),( 6, 9)), 1, 10) -- 13534
,( 11, E,0,0,((46,49),(35,35),( 6, 7),(20,20),(16,17),( 8,11)), 1, 10) -- 13535
,( 11, E,0,0,((38,41),(28,29),( 0, 1),(14,15),(14,15),(10,13)), 1, 10) -- 13536
,( 11, E,0,0,((40,43),(30,31),( 2, 3),(16,17),(16,17),(12,15)), 1, 10) -- 13537
,( 11, E,0,0,((42,45),(32,33),( 4, 5),(18,19),(18,19),(14,17)), 1, 10) -- 13538
,( 11, E,0,0,((44,47),(34,35),( 6, 7),(20,21),(20,21),(16,19)), 1, 10) -- 13539
,( 11, E,0,0,((42,42),(29,29),( 0, 0),(13,13),(10,10),( 0, 3)), 1, 10) -- 13540
,( 11, E,0,0,((44,44),(31,31),( 2, 2),(15,15),(12,12),( 2, 5)), 1, 10) -- 13541
,( 11, E,0,0,((46,46),(33,33),( 4, 4),(17,17),(14,14),( 4, 7)), 1, 10) -- 13542
,( 11, E,0,0,((48,48),(35,35),( 6, 6),(19,19),(16,16),( 6, 9)), 1, 10) -- 13543
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 4, 7)), 1,  9) -- 13544
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 6, 9)), 1,  9) -- 13545
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 8,11)), 1,  9) -- 13546
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(10,13)), 1,  9) -- 13547
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),( 8,11)), 1,  9) -- 13548
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),(10,13)), 1,  9) -- 13549
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),(12,15)), 1,  9) -- 13550
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(14,17)), 1,  9) -- 13551
,( 11, E,0,0,((40,43),(28,29),( 0, 0),(13,13),(12,13),( 8,11)), 1,  9) -- 13552
,( 11, E,0,0,((42,45),(30,31),( 2, 2),(15,15),(14,15),(10,13)), 1,  9) -- 13553
,( 11, E,0,0,((44,47),(32,33),( 4, 4),(17,17),(16,17),(12,15)), 1,  9) -- 13554
,( 11, E,0,0,((46,49),(34,35),( 6, 6),(19,19),(18,19),(14,17)), 1,  9) -- 13555
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 13556
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 13557
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 13558
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 13559
,( 11, E,0,0,((40,43),(29,29),( 0, 0),(12,13),(10,11),( 4, 7)), 1,  9) -- 13560
,( 11, E,0,0,((42,45),(31,31),( 2, 2),(14,15),(12,13),( 6, 9)), 1,  9) -- 13561
,( 11, E,0,0,((44,47),(33,33),( 4, 4),(16,17),(14,15),( 8,11)), 1,  9) -- 13562
,( 11, E,0,0,((46,49),(35,35),( 6, 6),(18,19),(16,17),(10,13)), 1,  9) -- 13563
,( 11, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(14,15),( 6, 9)), 1,  9) -- 13564
,( 11, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(16,17),( 8,11)), 1,  9) -- 13565
,( 11, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(18,19),(10,13)), 1,  9) -- 13566
,( 11, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(20,21),(12,15)), 1,  9) -- 13567
,( 11, E,0,0,((40,43),(29,29),( 0, 1),(14,14),(12,13),( 8,11)), 1,  9) -- 13568
,( 11, E,0,0,((42,45),(31,31),( 2, 3),(16,16),(14,15),(10,13)), 1,  9) -- 13569
,( 11, E,0,0,((44,47),(33,33),( 4, 5),(18,18),(16,17),(12,15)), 1,  9) -- 13570
,( 11, E,0,0,((46,49),(35,35),( 6, 7),(20,20),(18,19),(14,17)), 1,  9) -- 13571
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 0, 3)), 1,  9) -- 13572
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),( 2, 5)), 1,  9) -- 13573
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),( 4, 7)), 1,  9) -- 13574
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),( 6, 9)), 1,  9) -- 13575
,( 11, E,0,0,((40,43),(28,29),( 0, 1),(12,13),( 8, 9),( 0, 3)), 1,  9) -- 13576
,( 11, E,0,0,((42,45),(30,31),( 2, 3),(14,15),(10,11),( 2, 5)), 1,  9) -- 13577
,( 11, E,0,0,((44,47),(32,33),( 4, 5),(16,17),(12,13),( 4, 7)), 1,  9) -- 13578
,( 11, E,0,0,((46,49),(34,35),( 6, 7),(18,19),(14,15),( 6, 9)), 1,  9) -- 13579
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(12,13),(10,11),( 8, 9)), 1,  9) -- 13580
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(14,15),(12,13),(10,11)), 1,  9) -- 13581
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(16,17),(14,15),(12,13)), 1,  9) -- 13582
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(18,19),(16,17),(14,15)), 1,  9) -- 13583
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(14,15),(12,13),( 4, 7)), 1,  9) -- 13584
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(16,17),(14,15),( 6, 9)), 1,  9) -- 13585
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(18,19),(16,17),( 8,11)), 1,  9) -- 13586
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(20,21),(18,19),(10,13)), 1,  9) -- 13587
,( 11, E,0,0,((40,43),(30,31),( 1, 1),(14,15),(14,14),(10,13)), 1,  9) -- 13588
,( 11, E,0,0,((42,45),(32,33),( 3, 3),(16,17),(16,16),(12,15)), 1,  9) -- 13589
,( 11, E,0,0,((44,47),(34,35),( 5, 5),(18,19),(18,18),(14,17)), 1,  9) -- 13590
,( 11, E,0,0,((46,49),(36,37),( 7, 7),(20,21),(20,20),(16,19)), 1,  9) -- 13591
,( 11, E,0,0,((42,42),(29,29),( 0, 1),(14,14),(12,13),( 4, 7)), 1,  9) -- 13592
,( 11, E,0,0,((44,44),(31,31),( 2, 3),(16,16),(14,15),( 6, 9)), 1,  9) -- 13593
,( 11, E,0,0,((46,46),(33,33),( 4, 5),(18,18),(16,17),( 8,11)), 1,  9) -- 13594
,( 11, E,0,0,((48,48),(35,35),( 6, 7),(20,20),(18,19),(10,13)), 1,  9) -- 13595
,( 11, E,0,0,((42,45),(30,31),( 1, 1),(14,15),(10,11),( 6, 7)), 1,  9) -- 13596
,( 11, E,0,0,((44,47),(32,33),( 3, 3),(16,17),(12,13),( 8, 9)), 1,  9) -- 13597
,( 11, E,0,0,((46,49),(34,35),( 5, 5),(18,19),(14,15),(10,11)), 1,  9) -- 13598
,( 11, E,0,0,((48,51),(36,37),( 7, 7),(20,21),(16,17),(12,13)), 1,  9) -- 13599
,( 11, E,0,0,((42,45),(30,31),( 0, 1),(13,13),(12,12),(10,13)), 1,  9) -- 13600
,( 11, E,0,0,((44,47),(32,33),( 2, 3),(15,15),(14,14),(12,15)), 1,  9) -- 13601
,( 11, E,0,0,((46,49),(34,35),( 4, 5),(17,17),(16,16),(14,17)), 1,  9) -- 13602
,( 11, E,0,0,((48,51),(36,37),( 6, 7),(19,19),(18,18),(16,19)), 1,  9) -- 13603
,( 11, E,0,0,((40,43),(28,29),( 0, 1),(14,15),(14,15),(14,15)), 1,  9) -- 13604
,( 11, E,0,0,((42,45),(30,31),( 2, 3),(16,17),(16,17),(16,17)), 1,  9) -- 13605
,( 11, E,0,0,((44,47),(32,33),( 4, 5),(18,19),(18,19),(18,19)), 1,  9) -- 13606
,( 11, E,0,0,((46,49),(34,35),( 6, 7),(20,21),(20,21),(20,21)), 1,  9) -- 13607
,( 11, E,0,0,((44,47),(30,33),( 0, 1),(12,15),(10,13),(12,15)), 1,  8) -- 13608
,( 11, E,0,0,((46,49),(32,35),( 2, 3),(14,17),(12,15),(14,17)), 1,  8) -- 13609
,( 11, E,0,0,((48,51),(34,37),( 4, 5),(16,19),(14,17),(16,19)), 1,  8) -- 13610
,( 11, E,0,0,((50,53),(36,39),( 6, 7),(18,21),(16,19),(18,21)), 1,  8) -- 13611
,( 11, E,0,0,((44,47),(30,33),( 0, 1),(10,13),( 6, 9),( 2, 5)), 1,  8) -- 13612
,( 11, E,0,0,((46,49),(32,35),( 2, 3),(12,15),( 8,11),( 4, 7)), 1,  8) -- 13613
,( 11, E,0,0,((48,51),(34,37),( 4, 5),(14,17),(10,13),( 6, 9)), 1,  8) -- 13614
,( 11, E,0,0,((50,53),(36,39),( 6, 7),(16,19),(12,15),( 8,11)), 1,  8) -- 13615
,( 11, E,0,0,((42,45),(28,31),( 0, 1),(12,15),(14,17),(14,14)), 1,  8) -- 13616
,( 11, E,0,0,((44,47),(30,33),( 2, 3),(14,17),(16,19),(16,16)), 1,  8) -- 13617
,( 11, E,0,0,((46,49),(32,35),( 4, 5),(16,19),(18,21),(18,18)), 1,  8) -- 13618
,( 11, E,0,0,((48,51),(34,37),( 6, 7),(18,21),(20,23),(20,20)), 1,  8) -- 13619
,( 11, E,0,0,((40,43),(28,31),( 0, 1),(12,15),(12,15),(10,13)), 1,  8) -- 13620
,( 11, E,0,0,((42,45),(30,33),( 2, 3),(14,17),(14,17),(12,15)), 1,  8) -- 13621
,( 11, E,0,0,((44,47),(32,35),( 4, 5),(16,19),(16,19),(14,17)), 1,  8) -- 13622
,( 11, E,0,0,((46,49),(34,37),( 6, 7),(18,21),(18,21),(16,19)), 1,  8) -- 13623
,( 11, E,0,0,((46,49),(30,33),( 0, 1),(10,13),(10,13),(99,99)), 1,  7) -- 13624
,( 11, E,0,0,((48,51),(32,35),( 2, 3),(12,15),(12,15),(99,99)), 1,  7) -- 13625
,( 11, E,0,0,((50,53),(34,37),( 4, 5),(14,17),(14,17),(99,99)), 1,  7) -- 13626
,( 11, E,0,0,((52,55),(36,39),( 6, 7),(16,19),(16,19),(99,99)), 1,  7) -- 13627
,( 11, E,0,0,((46,49),(30,33),( 0, 1),(12,15),(14,17),(99,99)), 1,  7) -- 13628
,( 11, E,0,0,((48,51),(32,35),( 2, 3),(14,17),(16,19),(99,99)), 1,  7) -- 13629
,( 11, E,0,0,((50,53),(34,37),( 4, 5),(16,19),(18,21),(99,99)), 1,  7) -- 13630
,( 11, E,0,0,((52,55),(36,39),( 6, 7),(18,21),(20,23),(99,99)), 1,  7) -- 13631
,( 11, E,0,1,((48,51),(32,35),( 0, 1),(10,13),(99,99),(99,99)), 1,  7) -- 13632
,( 11, E,0,1,((50,53),(34,37),( 2, 3),(12,15),(99,99),(99,99)), 1,  7) -- 13633
,( 11, E,0,1,((52,55),(36,39),( 4, 5),(14,17),(99,99),(99,99)), 1,  7) -- 13634
,( 11, E,0,1,((54,57),(38,41),( 6, 7),(16,19),(99,99),(99,99)), 1,  7) -- 13635
,( 11, E,0,1,((46,49),(30,33),( 0, 1),(14,17),(99,99),(99,99)), 1,  7) -- 13636
,( 11, E,0,1,((48,51),(32,35),( 2, 3),(16,19),(99,99),(99,99)), 1,  7) -- 13637
,( 11, E,0,1,((50,53),(34,37),( 4, 5),(18,21),(99,99),(99,99)), 1,  7) -- 13638
,( 11, E,0,1,((52,55),(36,39),( 6, 7),(20,23),(99,99),(99,99)), 1,  7) -- 13639
,( 11, E,0,1,((50,53),(32,35),( 0, 1),(12,15),(99,99),(99,99)), 1,  6) -- 13640
,( 11, E,0,1,((52,55),(34,37),( 2, 3),(14,17),(99,99),(99,99)), 1,  6) -- 13641
,( 11, E,0,1,((54,57),(36,39),( 4, 5),(16,19),(99,99),(99,99)), 1,  6) -- 13642
,( 11, E,0,1,((56,59),(38,41),( 6, 7),(18,21),(99,99),(99,99)), 1,  6) -- 13643
,( 11, E,0,1,((42,45),(28,31),( 0, 1),(16,19),(99,99),(99,99)), 1,  6) -- 13644
,( 11, E,0,1,((44,47),(30,33),( 2, 3),(18,21),(99,99),(99,99)), 1,  6) -- 13645
,( 11, E,0,1,((46,49),(32,35),( 4, 5),(20,23),(99,99),(99,99)), 1,  6) -- 13646
,( 11, E,0,1,((48,51),(34,37),( 6, 7),(22,25),(99,99),(99,99)), 1,  6) -- 13647
,( 11, E,0,1,((40,43),(26,29),( 0, 1),(16,17),(99,99),(99,99)), 1,  5) -- 13648
,( 11, E,0,1,((42,45),(28,31),( 2, 3),(18,19),(99,99),(99,99)), 1,  5) -- 13649
,( 11, E,0,1,((44,47),(30,33),( 4, 5),(20,21),(99,99),(99,99)), 1,  5) -- 13650
,( 11, E,0,1,((46,49),(32,35),( 6, 7),(22,23),(99,99),(99,99)), 1,  5) -- 13651
,( 11, E,0,1,((54,57),(36,37),( 0, 1),(12,13),(99,99),(99,99)), 1,  5) -- 13652
,( 11, E,0,1,((56,59),(38,39),( 2, 3),(14,15),(99,99),(99,99)), 1,  5) -- 13653
,( 11, E,0,1,((58,61),(40,41),( 4, 5),(16,17),(99,99),(99,99)), 1,  5) -- 13654
,( 11, E,0,1,((60,63),(42,43),( 6, 7),(18,19),(99,99),(99,99)), 1,  5) -- 13655
,( 11, E,0,1,((46,47),(30,31),( 0, 1),(18,19),(99,99),(99,99)), 1,  5) -- 13656
,( 11, E,0,1,((48,49),(32,33),( 2, 3),(20,21),(99,99),(99,99)), 1,  5) -- 13657
,( 11, E,0,1,((50,51),(34,35),( 4, 5),(22,23),(99,99),(99,99)), 1,  5) -- 13658
,( 11, E,0,1,((52,53),(36,37),( 6, 7),(24,25),(99,99),(99,99)), 1,  5) -- 13659
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 13660
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 13661
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 13662
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 13663
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 13664
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 13665
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 13666
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 13667
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 13668
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 13669
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 13670
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 13671
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 13672
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 13673
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 13674
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 13675
,( 11, E,0,0,((31,31),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 31) -- 13676
,( 11, E,0,0,((32,32),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 31) -- 13677
,( 11, E,0,0,((33,33),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 31) -- 13678
,( 11, E,0,0,((34,34),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 31) -- 13679
,( 11, E,0,0,((35,35),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 31) -- 13680
,( 11, E,0,0,((36,36),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 31) -- 13681
,( 11, E,0,0,((37,37),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 31) -- 13682
,( 11, E,0,0,((38,38),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 31) -- 13683
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 31) -- 13684
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 31) -- 13685
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(10,10)), 0, 31) -- 13686
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(11,11)), 0, 31) -- 13687
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(12,12)), 0, 31) -- 13688
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(13,13)), 0, 31) -- 13689
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(14,14)), 0, 31) -- 13690
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(15,15)), 0, 31) -- 13691
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 31) -- 13692
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 31) -- 13693
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 31) -- 13694
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 31) -- 13695
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 31) -- 13696
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 31) -- 13697
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 31) -- 13698
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 31) -- 13699
,( 11, E,0,0,((32,32),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 31) -- 13700
,( 11, E,0,0,((33,33),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 31) -- 13701
,( 11, E,0,0,((34,34),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 31) -- 13702
,( 11, E,0,0,((35,35),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 31) -- 13703
,( 11, E,0,0,((36,36),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 31) -- 13704
,( 11, E,0,0,((37,37),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 31) -- 13705
,( 11, E,0,0,((38,38),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 31) -- 13706
,( 11, E,0,0,((39,39),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 31) -- 13707
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 30) -- 13708
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(17,17),(10,10)), 0, 30) -- 13709
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(18,18),(11,11)), 0, 30) -- 13710
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(19,19),(12,12)), 0, 30) -- 13711
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(20,20),(13,13)), 0, 30) -- 13712
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(21,21),(14,14)), 0, 30) -- 13713
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(22,22),(15,15)), 0, 30) -- 13714
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(23,23),(16,16)), 0, 30) -- 13715
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 28) -- 13716
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(10,10)), 0, 28) -- 13717
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(11,11)), 0, 28) -- 13718
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(12,12)), 0, 28) -- 13719
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(13,13)), 0, 28) -- 13720
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(14,14)), 0, 28) -- 13721
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(15,15)), 0, 28) -- 13722
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(16,16)), 0, 28) -- 13723
,( 11, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 27) -- 13724
,( 11, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 27) -- 13725
,( 11, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 27) -- 13726
,( 11, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 27) -- 13727
,( 11, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 27) -- 13728
,( 11, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 27) -- 13729
,( 11, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 27) -- 13730
,( 11, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 27) -- 13731
,( 11, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 26) -- 13732
,( 11, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 26) -- 13733
,( 11, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 26) -- 13734
,( 11, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 26) -- 13735
,( 11, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 26) -- 13736
,( 11, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 26) -- 13737
,( 11, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 26) -- 13738
,( 11, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 26) -- 13739
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 8, 8)), 0, 24) -- 13740
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),( 9, 9)), 0, 24) -- 13741
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(10,10)), 0, 24) -- 13742
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(11,11)), 0, 24) -- 13743
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(12,12)), 0, 24) -- 13744
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(13,13)), 0, 24) -- 13745
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(14,14)), 0, 24) -- 13746
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(15,15)), 0, 24) -- 13747
,( 11, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 24) -- 13748
,( 11, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 24) -- 13749
,( 11, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 24) -- 13750
,( 11, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 24) -- 13751
,( 11, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 24) -- 13752
,( 11, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 24) -- 13753
,( 11, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 24) -- 13754
,( 11, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 24) -- 13755
,( 11, E,0,0,((31,31),(24,24),( 0, 0),(16,16),(17,17),(10,10)), 0, 24) -- 13756
,( 11, E,0,0,((32,32),(25,25),( 1, 1),(17,17),(18,18),(11,11)), 0, 24) -- 13757
,( 11, E,0,0,((33,33),(26,26),( 2, 2),(18,18),(19,19),(12,12)), 0, 24) -- 13758
,( 11, E,0,0,((34,34),(27,27),( 3, 3),(19,19),(20,20),(13,13)), 0, 24) -- 13759
,( 11, E,0,0,((35,35),(28,28),( 4, 4),(20,20),(21,21),(14,14)), 0, 24) -- 13760
,( 11, E,0,0,((36,36),(29,29),( 5, 5),(21,21),(22,22),(15,15)), 0, 24) -- 13761
,( 11, E,0,0,((37,37),(30,30),( 6, 6),(22,22),(23,23),(16,16)), 0, 24) -- 13762
,( 11, E,0,0,((38,38),(31,31),( 7, 7),(23,23),(24,24),(17,17)), 0, 24) -- 13763
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 9, 9)), 0, 23) -- 13764
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),(10,10)), 0, 23) -- 13765
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(11,11)), 0, 23) -- 13766
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(12,12)), 0, 23) -- 13767
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(13,13)), 0, 23) -- 13768
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(14,14)), 0, 23) -- 13769
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(15,15)), 0, 23) -- 13770
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(16,16)), 0, 23) -- 13771
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(15,15),(16,16),( 9, 9)), 0, 23) -- 13772
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(16,16),(17,17),(10,10)), 0, 23) -- 13773
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(17,17),(18,18),(11,11)), 0, 23) -- 13774
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(18,18),(19,19),(12,12)), 0, 23) -- 13775
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(19,19),(20,20),(13,13)), 0, 23) -- 13776
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(20,20),(21,21),(14,14)), 0, 23) -- 13777
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(21,21),(22,22),(15,15)), 0, 23) -- 13778
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(22,22),(23,23),(16,16)), 0, 23) -- 13779
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 22) -- 13780
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 22) -- 13781
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 22) -- 13782
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 22) -- 13783
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 22) -- 13784
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 22) -- 13785
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 22) -- 13786
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 22) -- 13787
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 21) -- 13788
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 21) -- 13789
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 21) -- 13790
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 21) -- 13791
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 21) -- 13792
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 21) -- 13793
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 21) -- 13794
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 21) -- 13795
,( 11, E,0,0,((31,31),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 20) -- 13796
,( 11, E,0,0,((32,32),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 20) -- 13797
,( 11, E,0,0,((33,33),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 20) -- 13798
,( 11, E,0,0,((34,34),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 20) -- 13799
,( 11, E,0,0,((35,35),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 20) -- 13800
,( 11, E,0,0,((36,36),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 20) -- 13801
,( 11, E,0,0,((37,37),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 20) -- 13802
,( 11, E,0,0,((38,38),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 20) -- 13803
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 19) -- 13804
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 19) -- 13805
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 19) -- 13806
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 19) -- 13807
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 19) -- 13808
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 19) -- 13809
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 19) -- 13810
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 19) -- 13811
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 19) -- 13812
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 19) -- 13813
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 19) -- 13814
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 19) -- 13815
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 19) -- 13816
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 19) -- 13817
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 19) -- 13818
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 19) -- 13819
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),(10,10)), 0, 19) -- 13820
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(11,11)), 0, 19) -- 13821
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(12,12)), 0, 19) -- 13822
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(13,13)), 0, 19) -- 13823
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(14,14)), 0, 19) -- 13824
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(15,15)), 0, 19) -- 13825
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(16,16)), 0, 19) -- 13826
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(17,17)), 0, 19) -- 13827
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 19) -- 13828
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(18,18),(10,10)), 0, 19) -- 13829
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(19,19),(11,11)), 0, 19) -- 13830
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(20,20),(12,12)), 0, 19) -- 13831
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(21,21),(13,13)), 0, 19) -- 13832
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(22,22),(14,14)), 0, 19) -- 13833
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(23,23),(15,15)), 0, 19) -- 13834
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(24,24),(16,16)), 0, 19) -- 13835
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(16,16),(16,16),( 8, 8)), 0, 19) -- 13836
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(17,17),(17,17),( 9, 9)), 0, 19) -- 13837
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(18,18),(18,18),(10,10)), 0, 19) -- 13838
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(19,19),(19,19),(11,11)), 0, 19) -- 13839
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(20,20),(20,20),(12,12)), 0, 19) -- 13840
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(21,21),(21,21),(13,13)), 0, 19) -- 13841
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(22,22),(22,22),(14,14)), 0, 19) -- 13842
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(23,23),(23,23),(15,15)), 0, 19) -- 13843
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 18) -- 13844
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 18) -- 13845
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 18) -- 13846
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 18) -- 13847
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 18) -- 13848
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 18) -- 13849
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 18) -- 13850
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 18) -- 13851
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 18) -- 13852
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 18) -- 13853
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 18) -- 13854
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 18) -- 13855
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 18) -- 13856
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 18) -- 13857
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 18) -- 13858
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 18) -- 13859
,( 11, E,0,0,((30,30),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 18) -- 13860
,( 11, E,0,0,((31,31),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 18) -- 13861
,( 11, E,0,0,((32,32),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 18) -- 13862
,( 11, E,0,0,((33,33),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 18) -- 13863
,( 11, E,0,0,((34,34),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 18) -- 13864
,( 11, E,0,0,((35,35),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 18) -- 13865
,( 11, E,0,0,((36,36),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 18) -- 13866
,( 11, E,0,0,((37,37),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 18) -- 13867
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(10,10)), 0, 18) -- 13868
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(11,11)), 0, 18) -- 13869
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(12,12)), 0, 18) -- 13870
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(13,13)), 0, 18) -- 13871
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(14,14)), 0, 18) -- 13872
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(15,15)), 0, 18) -- 13873
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(16,16)), 0, 18) -- 13874
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(17,17)), 0, 18) -- 13875
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(11,11)), 0, 17) -- 13876
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(12,12)), 0, 17) -- 13877
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(13,13)), 0, 17) -- 13878
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(14,14)), 0, 17) -- 13879
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(15,15)), 0, 17) -- 13880
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(16,16)), 0, 17) -- 13881
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(17,17)), 0, 17) -- 13882
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(18,18)), 0, 17) -- 13883
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 17) -- 13884
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 17) -- 13885
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 17) -- 13886
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 17) -- 13887
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 17) -- 13888
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 17) -- 13889
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 17) -- 13890
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 17) -- 13891
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(16,16),(18,18),(11,11)), 0, 17) -- 13892
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(17,17),(19,19),(12,12)), 0, 17) -- 13893
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(18,18),(20,20),(13,13)), 0, 17) -- 13894
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(19,19),(21,21),(14,14)), 0, 17) -- 13895
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(20,20),(22,22),(15,15)), 0, 17) -- 13896
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(21,21),(23,23),(16,16)), 0, 17) -- 13897
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(22,22),(24,24),(17,17)), 0, 17) -- 13898
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(23,23),(25,25),(18,18)), 0, 17) -- 13899
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(18,18),(10,10)), 0, 17) -- 13900
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(19,19),(11,11)), 0, 17) -- 13901
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(20,20),(12,12)), 0, 17) -- 13902
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(21,21),(13,13)), 0, 17) -- 13903
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(22,22),(14,14)), 0, 17) -- 13904
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(23,23),(15,15)), 0, 17) -- 13905
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(24,24),(16,16)), 0, 17) -- 13906
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(25,25),(17,17)), 0, 17) -- 13907
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 13908
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 13909
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 13910
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 13911
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 13912
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 13913
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 13914
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 13915
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(16,16),(18,18),(11,11)), 0, 16) -- 13916
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(17,17),(19,19),(12,12)), 0, 16) -- 13917
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(18,18),(20,20),(13,13)), 0, 16) -- 13918
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(19,19),(21,21),(14,14)), 0, 16) -- 13919
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(20,20),(22,22),(15,15)), 0, 16) -- 13920
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(21,21),(23,23),(16,16)), 0, 16) -- 13921
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(22,22),(24,24),(17,17)), 0, 16) -- 13922
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(23,23),(25,25),(18,18)), 0, 16) -- 13923
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(18,18),(10,10)), 0, 16) -- 13924
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(19,19),(11,11)), 0, 16) -- 13925
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(20,20),(12,12)), 0, 16) -- 13926
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(21,21),(13,13)), 0, 16) -- 13927
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(22,22),(14,14)), 0, 16) -- 13928
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(23,23),(15,15)), 0, 16) -- 13929
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(24,24),(16,16)), 0, 16) -- 13930
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(25,25),(17,17)), 0, 16) -- 13931
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),(10,10)), 0, 16) -- 13932
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(11,11)), 0, 16) -- 13933
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(12,12)), 0, 16) -- 13934
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(13,13)), 0, 16) -- 13935
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(14,14)), 0, 16) -- 13936
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(15,15)), 0, 16) -- 13937
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(16,16)), 0, 16) -- 13938
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(17,17)), 0, 16) -- 13939
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(12,12)), 0, 16) -- 13940
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(13,13)), 0, 16) -- 13941
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(14,14)), 0, 16) -- 13942
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(15,15)), 0, 16) -- 13943
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(16,16)), 0, 16) -- 13944
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(17,17)), 0, 16) -- 13945
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(18,18)), 0, 16) -- 13946
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(19,19)), 0, 16) -- 13947
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 13948
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 13949
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 13950
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 13951
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 13952
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 13953
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 13954
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 13955
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(18,18),(11,11)), 0, 15) -- 13956
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(19,19),(12,12)), 0, 15) -- 13957
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(20,20),(13,13)), 0, 15) -- 13958
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(21,21),(14,14)), 0, 15) -- 13959
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(22,22),(15,15)), 0, 15) -- 13960
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(23,23),(16,16)), 0, 15) -- 13961
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(24,24),(17,17)), 0, 15) -- 13962
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(25,25),(18,18)), 0, 15) -- 13963
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(17,17),(19,19),(12,12)), 0, 15) -- 13964
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(18,18),(20,20),(13,13)), 0, 15) -- 13965
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(19,19),(21,21),(14,14)), 0, 15) -- 13966
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(20,20),(22,22),(15,15)), 0, 15) -- 13967
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(21,21),(23,23),(16,16)), 0, 15) -- 13968
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(22,22),(24,24),(17,17)), 0, 15) -- 13969
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(23,23),(25,25),(18,18)), 0, 15) -- 13970
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(24,24),(26,26),(19,19)), 0, 15) -- 13971
,( 11, E,0,0,((29,29),(23,23),( 0, 0),(17,17),(19,19),(11,11)), 0, 15) -- 13972
,( 11, E,0,0,((30,30),(24,24),( 1, 1),(18,18),(20,20),(12,12)), 0, 15) -- 13973
,( 11, E,0,0,((31,31),(25,25),( 2, 2),(19,19),(21,21),(13,13)), 0, 15) -- 13974
,( 11, E,0,0,((32,32),(26,26),( 3, 3),(20,20),(22,22),(14,14)), 0, 15) -- 13975
,( 11, E,0,0,((33,33),(27,27),( 4, 4),(21,21),(23,23),(15,15)), 0, 15) -- 13976
,( 11, E,0,0,((34,34),(28,28),( 5, 5),(22,22),(24,24),(16,16)), 0, 15) -- 13977
,( 11, E,0,0,((35,35),(29,29),( 6, 6),(23,23),(25,25),(17,17)), 0, 15) -- 13978
,( 11, E,0,0,((36,36),(30,30),( 7, 7),(24,24),(26,26),(18,18)), 0, 15) -- 13979
,( 11, E,0,0,((28,28),(22,22),( 0, 0),(16,16),(17,17),( 9, 9)), 0, 15) -- 13980
,( 11, E,0,0,((29,29),(23,23),( 1, 1),(17,17),(18,18),(10,10)), 0, 15) -- 13981
,( 11, E,0,0,((30,30),(24,24),( 2, 2),(18,18),(19,19),(11,11)), 0, 15) -- 13982
,( 11, E,0,0,((31,31),(25,25),( 3, 3),(19,19),(20,20),(12,12)), 0, 15) -- 13983
,( 11, E,0,0,((32,32),(26,26),( 4, 4),(20,20),(21,21),(13,13)), 0, 15) -- 13984
,( 11, E,0,0,((33,33),(27,27),( 5, 5),(21,21),(22,22),(14,14)), 0, 15) -- 13985
,( 11, E,0,0,((34,34),(28,28),( 6, 6),(22,22),(23,23),(15,15)), 0, 15) -- 13986
,( 11, E,0,0,((35,35),(29,29),( 7, 7),(23,23),(24,24),(16,16)), 0, 15) -- 13987
,( 11, E,0,0,((29,29),(22,22),( 0, 0),(17,17),(18,18),(10,10)), 0, 15) -- 13988
,( 11, E,0,0,((30,30),(23,23),( 1, 1),(18,18),(19,19),(11,11)), 0, 15) -- 13989
,( 11, E,0,0,((31,31),(24,24),( 2, 2),(19,19),(20,20),(12,12)), 0, 15) -- 13990
,( 11, E,0,0,((32,32),(25,25),( 3, 3),(20,20),(21,21),(13,13)), 0, 15) -- 13991
,( 11, E,0,0,((33,33),(26,26),( 4, 4),(21,21),(22,22),(14,14)), 0, 15) -- 13992
,( 11, E,0,0,((34,34),(27,27),( 5, 5),(22,22),(23,23),(15,15)), 0, 15) -- 13993
,( 11, E,0,0,((35,35),(28,28),( 6, 6),(23,23),(24,24),(16,16)), 0, 15) -- 13994
,( 11, E,0,0,((36,36),(29,29),( 7, 7),(24,24),(25,25),(17,17)), 0, 15) -- 13995
,( 11, E,0,0,((26,29),(22,23),( 0, 1),(16,17),(18,19),(10,13)), 0, 14) -- 13996
,( 11, E,0,0,((28,31),(24,25),( 2, 3),(18,19),(20,21),(12,15)), 0, 14) -- 13997
,( 11, E,0,0,((30,33),(26,27),( 4, 5),(20,21),(22,23),(14,17)), 0, 14) -- 13998
,( 11, E,0,0,((32,35),(28,29),( 6, 7),(22,23),(24,25),(16,19)), 0, 14) -- 13999
,( 11, E,0,0,((28,31),(22,23),( 1, 1),(18,18),(20,21),(12,15)), 0, 14) -- 14000
,( 11, E,0,0,((30,33),(24,25),( 3, 3),(20,20),(22,23),(14,17)), 0, 14) -- 14001
,( 11, E,0,0,((32,35),(26,27),( 5, 5),(22,22),(24,25),(16,19)), 0, 14) -- 14002
,( 11, E,0,0,((34,37),(28,29),( 7, 7),(24,24),(26,27),(18,21)), 0, 14) -- 14003
,( 11, E,0,0,((26,29),(21,21),( 0, 0),(16,17),(18,19),(10,13)), 0, 14) -- 14004
,( 11, E,0,0,((28,31),(23,23),( 2, 2),(18,19),(20,21),(12,15)), 0, 14) -- 14005
,( 11, E,0,0,((30,33),(25,25),( 4, 4),(20,21),(22,23),(14,17)), 0, 14) -- 14006
,( 11, E,0,0,((32,35),(27,27),( 6, 6),(22,23),(24,25),(16,19)), 0, 14) -- 14007
,( 11, E,0,0,((26,29),(22,23),( 0, 1),(18,18),(19,19),(10,13)), 0, 13) -- 14008
,( 11, E,0,0,((28,31),(24,25),( 2, 3),(20,20),(21,21),(12,15)), 0, 13) -- 14009
,( 11, E,0,0,((30,33),(26,27),( 4, 5),(22,22),(23,23),(14,17)), 0, 13) -- 14010
,( 11, E,0,0,((32,35),(28,29),( 6, 7),(24,24),(25,25),(16,19)), 0, 13) -- 14011
,( 11, E,0,0,((26,29),(22,23),( 0, 1),(18,19),(20,21),(12,15)), 0, 13) -- 14012
,( 11, E,0,0,((28,31),(24,25),( 2, 3),(20,21),(22,23),(14,17)), 0, 13) -- 14013
,( 11, E,0,0,((30,33),(26,27),( 4, 5),(22,23),(24,25),(16,19)), 0, 13) -- 14014
,( 11, E,0,0,((32,35),(28,29),( 6, 7),(24,25),(26,27),(18,21)), 0, 13) -- 14015
,( 11, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(12,15)), 0, 12) -- 14016
,( 11, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(14,17)), 0, 12) -- 14017
,( 11, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(16,19)), 0, 12) -- 14018
,( 11, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(18,21)), 0, 12) -- 14019
,( 11, E,0,0,((24,27),(20,21),( 0, 0),(17,17),(20,21),(12,15)), 0, 12) -- 14020
,( 11, E,0,0,((26,29),(22,23),( 2, 2),(19,19),(22,23),(14,17)), 0, 12) -- 14021
,( 11, E,0,0,((28,31),(24,25),( 4, 4),(21,21),(24,25),(16,19)), 0, 12) -- 14022
,( 11, E,0,0,((30,33),(26,27),( 6, 6),(23,23),(26,27),(18,21)), 0, 12) -- 14023
,( 11, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(20,20),(10,11)), 0, 12) -- 14024
,( 11, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(22,22),(12,13)), 0, 12) -- 14025
,( 11, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(24,24),(14,15)), 0, 12) -- 14026
,( 11, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(26,26),(16,17)), 0, 12) -- 14027
,( 11, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(22,23),(14,17)), 0, 11) -- 14028
,( 11, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(24,25),(16,19)), 0, 11) -- 14029
,( 11, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(26,27),(18,21)), 0, 11) -- 14030
,( 11, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(28,29),(20,23)), 0, 11) -- 14031
,( 11, E,0,0,((24,27),(20,21),( 0, 0),(16,17),(18,19),( 8,11)), 0, 11) -- 14032
,( 11, E,0,0,((26,29),(22,23),( 2, 2),(18,19),(20,21),(10,13)), 0, 11) -- 14033
,( 11, E,0,0,((28,31),(24,25),( 4, 4),(20,21),(22,23),(12,15)), 0, 11) -- 14034
,( 11, E,0,0,((30,33),(26,27),( 6, 6),(22,23),(24,25),(14,17)), 0, 11) -- 14035
,( 11, E,0,0,((24,27),(20,21),( 0, 1),(18,19),(20,21),(10,11)), 0, 11) -- 14036
,( 11, E,0,0,((26,29),(22,23),( 2, 3),(20,21),(22,23),(12,13)), 0, 11) -- 14037
,( 11, E,0,0,((28,31),(24,25),( 4, 5),(22,23),(24,25),(14,15)), 0, 11) -- 14038
,( 11, E,0,0,((30,33),(26,27),( 6, 7),(24,25),(26,27),(16,17)), 0, 11) -- 14039
,( 11, E,0,0,((26,29),(22,23),( 1, 1),(18,19),(22,23),(14,17)), 0, 11) -- 14040
,( 11, E,0,0,((28,31),(24,25),( 3, 3),(20,21),(24,25),(16,19)), 0, 11) -- 14041
,( 11, E,0,0,((30,33),(26,27),( 5, 5),(22,23),(26,27),(18,21)), 0, 11) -- 14042
,( 11, E,0,0,((32,35),(28,29),( 7, 7),(24,25),(28,29),(20,23)), 0, 11) -- 14043
,( 11, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(20,20),(10,13)), 0, 11) -- 14044
,( 11, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(22,22),(12,15)), 0, 11) -- 14045
,( 11, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(24,24),(14,17)), 0, 11) -- 14046
,( 11, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(26,26),(16,19)), 0, 11) -- 14047
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),(12,15)), 0, 11) -- 14048
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(14,17)), 0, 11) -- 14049
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(16,19)), 0, 11) -- 14050
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(18,21)), 0, 11) -- 14051
,( 11, E,0,0,((24,27),(21,21),( 0, 1),(18,18),(19,19),(10,11)), 0, 11) -- 14052
,( 11, E,0,0,((26,29),(23,23),( 2, 3),(20,20),(21,21),(12,13)), 0, 11) -- 14053
,( 11, E,0,0,((28,31),(25,25),( 4, 5),(22,22),(23,23),(14,15)), 0, 11) -- 14054
,( 11, E,0,0,((30,33),(27,27),( 6, 7),(24,24),(25,25),(16,17)), 0, 11) -- 14055
,( 11, E,0,0,((20,23),(18,19),( 0, 0),(18,19),(20,21),(10,13)), 0, 10) -- 14056
,( 11, E,0,0,((22,25),(20,21),( 2, 2),(20,21),(22,23),(12,15)), 0, 10) -- 14057
,( 11, E,0,0,((24,27),(22,23),( 4, 4),(22,23),(24,25),(14,17)), 0, 10) -- 14058
,( 11, E,0,0,((26,29),(24,25),( 6, 6),(24,25),(26,27),(16,19)), 0, 10) -- 14059
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(12,15)), 0, 10) -- 14060
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(14,17)), 0, 10) -- 14061
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(16,19)), 0, 10) -- 14062
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(18,21)), 0, 10) -- 14063
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 8,11)), 0, 10) -- 14064
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),(10,13)), 0, 10) -- 14065
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),(12,15)), 0, 10) -- 14066
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(14,17)), 0, 10) -- 14067
,( 11, E,0,0,((23,23),(20,20),( 0, 1),(18,19),(20,21),(12,15)), 0, 10) -- 14068
,( 11, E,0,0,((25,25),(22,22),( 2, 3),(20,21),(22,23),(14,17)), 0, 10) -- 14069
,( 11, E,0,0,((27,27),(24,24),( 4, 5),(22,23),(24,25),(16,19)), 0, 10) -- 14070
,( 11, E,0,0,((29,29),(26,26),( 6, 7),(24,25),(26,27),(18,21)), 0, 10) -- 14071
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,18),(18,19),( 6, 9)), 0, 10) -- 14072
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,20),(20,21),( 8,11)), 0, 10) -- 14073
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,22),(22,23),(10,13)), 0, 10) -- 14074
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,24),(24,25),(12,15)), 0, 10) -- 14075
,( 11, E,0,0,((22,23),(19,19),( 0, 0),(18,18),(21,21),(14,17)), 0, 10) -- 14076
,( 11, E,0,0,((24,25),(21,21),( 2, 2),(20,20),(23,23),(16,19)), 0, 10) -- 14077
,( 11, E,0,0,((26,27),(23,23),( 4, 4),(22,22),(25,25),(18,21)), 0, 10) -- 14078
,( 11, E,0,0,((28,29),(25,25),( 6, 6),(24,24),(27,27),(20,23)), 0, 10) -- 14079
,( 11, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(14,17)), 0, 10) -- 14080
,( 11, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(16,19)), 0, 10) -- 14081
,( 11, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(18,21)), 0, 10) -- 14082
,( 11, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(20,23)), 0, 10) -- 14083
,( 11, E,0,0,((23,23),(19,19),( 0, 0),(17,17),(20,21),(10,13)), 0, 10) -- 14084
,( 11, E,0,0,((25,25),(21,21),( 2, 2),(19,19),(22,23),(12,15)), 0, 10) -- 14085
,( 11, E,0,0,((27,27),(23,23),( 4, 4),(21,21),(24,25),(14,17)), 0, 10) -- 14086
,( 11, E,0,0,((29,29),(25,25),( 6, 6),(23,23),(26,27),(16,19)), 0, 10) -- 14087
,( 11, E,0,0,((26,27),(22,22),( 1, 1),(18,19),(20,21),( 8,11)), 0, 10) -- 14088
,( 11, E,0,0,((28,29),(24,24),( 3, 3),(20,21),(22,23),(10,13)), 0, 10) -- 14089
,( 11, E,0,0,((30,31),(26,26),( 5, 5),(22,23),(24,25),(12,15)), 0, 10) -- 14090
,( 11, E,0,0,((32,33),(28,28),( 7, 7),(24,25),(26,27),(14,17)), 0, 10) -- 14091
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(17,17),(18,19),( 4, 7)), 0, 10) -- 14092
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(19,19),(20,21),( 6, 9)), 0, 10) -- 14093
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(21,21),(22,23),( 8,11)), 0, 10) -- 14094
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(23,23),(24,25),(10,13)), 0, 10) -- 14095
,( 11, E,0,0,((23,23),(20,20),( 0, 1),(19,19),(22,23),(16,17)), 0, 10) -- 14096
,( 11, E,0,0,((25,25),(22,22),( 2, 3),(21,21),(24,25),(18,19)), 0, 10) -- 14097
,( 11, E,0,0,((27,27),(24,24),( 4, 5),(23,23),(26,27),(20,21)), 0, 10) -- 14098
,( 11, E,0,0,((29,29),(26,26),( 6, 7),(25,25),(28,29),(22,23)), 0, 10) -- 14099
,( 11, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(24,25),(14,17)), 0, 10) -- 14100
,( 11, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(26,27),(16,19)), 0, 10) -- 14101
,( 11, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(28,29),(18,21)), 0, 10) -- 14102
,( 11, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(30,31),(20,23)), 0, 10) -- 14103
,( 11, E,0,0,((20,23),(19,19),( 0, 0),(18,19),(20,21),( 8, 9)), 0, 10) -- 14104
,( 11, E,0,0,((22,25),(21,21),( 2, 2),(20,21),(22,23),(10,11)), 0, 10) -- 14105
,( 11, E,0,0,((24,27),(23,23),( 4, 4),(22,23),(24,25),(12,13)), 0, 10) -- 14106
,( 11, E,0,0,((26,29),(25,25),( 6, 6),(24,25),(26,27),(14,15)), 0, 10) -- 14107
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(20,21),( 6, 9)), 0,  9) -- 14108
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(22,23),( 8,11)), 0,  9) -- 14109
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(24,25),(10,13)), 0,  9) -- 14110
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(26,27),(12,15)), 0,  9) -- 14111
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),( 8,11)), 0,  9) -- 14112
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(10,13)), 0,  9) -- 14113
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(12,15)), 0,  9) -- 14114
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(14,17)), 0,  9) -- 14115
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(20,21),(22,23),(10,13)), 0,  9) -- 14116
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(22,23),(24,25),(12,15)), 0,  9) -- 14117
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(24,25),(26,27),(14,17)), 0,  9) -- 14118
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(26,27),(28,29),(16,19)), 0,  9) -- 14119
,( 11, E,0,0,((22,25),(20,21),( 1, 1),(20,20),(22,23),(10,13)), 0,  9) -- 14120
,( 11, E,0,0,((24,27),(22,23),( 3, 3),(22,22),(24,25),(12,15)), 0,  9) -- 14121
,( 11, E,0,0,((26,29),(24,25),( 5, 5),(24,24),(26,27),(14,17)), 0,  9) -- 14122
,( 11, E,0,0,((28,31),(26,27),( 7, 7),(26,26),(28,29),(16,19)), 0,  9) -- 14123
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(20,21),( 4, 7)), 0,  9) -- 14124
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(22,23),( 6, 9)), 0,  9) -- 14125
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(24,25),( 8,11)), 0,  9) -- 14126
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(26,27),(10,13)), 0,  9) -- 14127
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(22,23),( 8,11)), 0,  9) -- 14128
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(24,25),(10,13)), 0,  9) -- 14129
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(26,27),(12,15)), 0,  9) -- 14130
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(28,29),(14,17)), 0,  9) -- 14131
,( 11, E,0,0,((18,21),(18,19),( 0, 1),(20,21),(24,25),(12,15)), 0,  9) -- 14132
,( 11, E,0,0,((20,23),(20,21),( 2, 3),(22,23),(26,27),(14,17)), 0,  9) -- 14133
,( 11, E,0,0,((22,25),(22,23),( 4, 5),(24,25),(28,29),(16,19)), 0,  9) -- 14134
,( 11, E,0,0,((24,27),(24,25),( 6, 7),(26,27),(30,31),(18,21)), 0,  9) -- 14135
,( 11, E,0,0,((22,25),(20,21),( 0, 1),(18,19),(18,19),( 2, 5)), 0,  9) -- 14136
,( 11, E,0,0,((24,27),(22,23),( 2, 3),(20,21),(20,21),( 4, 7)), 0,  9) -- 14137
,( 11, E,0,0,((26,29),(24,25),( 4, 5),(22,23),(22,23),( 6, 9)), 0,  9) -- 14138
,( 11, E,0,0,((28,31),(26,27),( 6, 7),(24,25),(24,25),( 8,11)), 0,  9) -- 14139
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(18,18),(18,19),( 4, 7)), 0,  9) -- 14140
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(20,20),(20,21),( 6, 9)), 0,  9) -- 14141
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(22,22),(22,23),( 8,11)), 0,  9) -- 14142
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(24,24),(24,25),(10,13)), 0,  9) -- 14143
,( 11, E,0,0,((18,21),(18,19),( 0, 1),(18,19),(20,21),( 4, 5)), 0,  9) -- 14144
,( 11, E,0,0,((20,23),(20,21),( 2, 3),(20,21),(22,23),( 6, 7)), 0,  9) -- 14145
,( 11, E,0,0,((22,25),(22,23),( 4, 5),(22,23),(24,25),( 8, 9)), 0,  9) -- 14146
,( 11, E,0,0,((24,27),(24,25),( 6, 7),(24,25),(26,27),(10,11)), 0,  9) -- 14147
,( 11, E,0,0,((18,21),(17,17),( 0, 0),(18,19),(22,23),(10,13)), 0,  9) -- 14148
,( 11, E,0,0,((20,23),(19,19),( 2, 2),(20,21),(24,25),(12,15)), 0,  9) -- 14149
,( 11, E,0,0,((22,25),(21,21),( 4, 4),(22,23),(26,27),(14,17)), 0,  9) -- 14150
,( 11, E,0,0,((24,27),(23,23),( 6, 6),(24,25),(28,29),(16,19)), 0,  9) -- 14151
,( 11, E,0,0,((20,23),(18,19),( 1, 1),(20,20),(24,25),(14,17)), 0,  9) -- 14152
,( 11, E,0,0,((22,25),(20,21),( 3, 3),(22,22),(26,27),(16,19)), 0,  9) -- 14153
,( 11, E,0,0,((24,27),(22,23),( 5, 5),(24,24),(28,29),(18,21)), 0,  9) -- 14154
,( 11, E,0,0,((26,29),(24,25),( 7, 7),(26,26),(30,31),(20,23)), 0,  9) -- 14155
,( 11, E,0,0,((20,23),(18,19),( 0, 0),(17,17),(18,19),( 6, 9)), 0,  9) -- 14156
,( 11, E,0,0,((22,25),(20,21),( 2, 2),(19,19),(20,21),( 8,11)), 0,  9) -- 14157
,( 11, E,0,0,((24,27),(22,23),( 4, 4),(21,21),(22,23),(10,13)), 0,  9) -- 14158
,( 11, E,0,0,((26,29),(24,25),( 6, 6),(23,23),(24,25),(12,15)), 0,  9) -- 14159
,( 11, E,0,0,((22,22),(19,19),( 1, 1),(19,19),(21,21),(10,13)), 0,  9) -- 14160
,( 11, E,0,0,((24,24),(21,21),( 3, 3),(21,21),(23,23),(12,15)), 0,  9) -- 14161
,( 11, E,0,0,((26,26),(23,23),( 5, 5),(23,23),(25,25),(14,17)), 0,  9) -- 14162
,( 11, E,0,0,((28,28),(25,25),( 7, 7),(25,25),(27,27),(16,19)), 0,  9) -- 14163
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(18,19),(22,23),(16,19)), 0,  9) -- 14164
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(20,21),(24,25),(18,21)), 0,  9) -- 14165
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(22,23),(26,27),(20,23)), 0,  9) -- 14166
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(24,25),(28,29),(22,23)), 0,  9) -- 14167
,( 11, E,0,0,((20,23),(20,20),( 1, 1),(20,20),(22,23),( 8,11)), 0,  9) -- 14168
,( 11, E,0,0,((22,25),(22,22),( 3, 3),(22,22),(24,25),(10,13)), 0,  9) -- 14169
,( 11, E,0,0,((24,27),(24,24),( 5, 5),(24,24),(26,27),(12,15)), 0,  9) -- 14170
,( 11, E,0,0,((26,29),(26,26),( 7, 7),(26,26),(28,29),(14,17)), 0,  9) -- 14171
,( 11, E,0,0,((16,19),(16,17),( 0, 0),(20,20),(24,25),(14,17)), 0,  9) -- 14172
,( 11, E,0,0,((18,21),(18,19),( 2, 2),(22,22),(26,27),(16,19)), 0,  9) -- 14173
,( 11, E,0,0,((20,23),(20,21),( 4, 4),(24,24),(28,29),(18,21)), 0,  9) -- 14174
,( 11, E,0,0,((22,25),(22,23),( 6, 6),(26,26),(30,31),(20,23)), 0,  9) -- 14175
,( 11, E,0,0,((18,21),(18,19),( 0, 1),(20,20),(22,23),(14,14)), 0,  9) -- 14176
,( 11, E,0,0,((20,23),(20,21),( 2, 3),(22,22),(24,25),(16,16)), 0,  9) -- 14177
,( 11, E,0,0,((22,25),(22,23),( 4, 5),(24,24),(26,27),(18,18)), 0,  9) -- 14178
,( 11, E,0,0,((24,27),(24,25),( 6, 7),(26,26),(28,29),(20,20)), 0,  9) -- 14179
,( 11, E,0,0,((18,21),(18,19),( 0, 1),(19,19),(22,22),( 6, 7)), 0,  9) -- 14180
,( 11, E,0,0,((20,23),(20,21),( 2, 3),(21,21),(24,24),( 8, 9)), 0,  9) -- 14181
,( 11, E,0,0,((22,25),(22,23),( 4, 5),(23,23),(26,26),(10,11)), 0,  9) -- 14182
,( 11, E,0,0,((24,27),(24,25),( 6, 7),(25,25),(28,28),(12,13)), 0,  9) -- 14183
,( 11, E,0,0,((22,25),(20,21),( 0, 0),(17,17),(16,17),( 5, 5)), 0,  9) -- 14184
,( 11, E,0,0,((24,27),(22,23),( 2, 2),(19,19),(18,19),( 7, 7)), 0,  9) -- 14185
,( 11, E,0,0,((26,29),(24,25),( 4, 4),(21,21),(20,21),( 9, 9)), 0,  9) -- 14186
,( 11, E,0,0,((28,31),(26,27),( 6, 6),(23,23),(22,23),(11,11)), 0,  9) -- 14187
,( 11, E,0,0,((18,21),(18,19),( 1, 1),(20,20),(23,23),( 8,11)), 0,  9) -- 14188
,( 11, E,0,0,((20,23),(20,21),( 3, 3),(22,22),(25,25),(10,13)), 0,  9) -- 14189
,( 11, E,0,0,((22,25),(22,23),( 5, 5),(24,24),(27,27),(12,15)), 0,  9) -- 14190
,( 11, E,0,0,((24,27),(24,25),( 7, 7),(26,26),(29,29),(14,17)), 0,  9) -- 14191
,( 11, E,0,0,((20,23),(18,19),( 0, 1),(19,19),(24,24),(14,17)), 0,  9) -- 14192
,( 11, E,0,0,((22,25),(20,21),( 2, 3),(21,21),(26,26),(16,19)), 0,  9) -- 14193
,( 11, E,0,0,((24,27),(22,23),( 4, 5),(23,23),(28,28),(18,21)), 0,  9) -- 14194
,( 11, E,0,0,((26,29),(24,25),( 6, 7),(25,25),(30,30),(20,23)), 0,  9) -- 14195
,( 11, E,0,0,((16,19),(17,17),( 0, 1),(18,19),(20,21),(99,99)), 0,  9) -- 14196
,( 11, E,0,0,((18,21),(19,19),( 2, 3),(20,21),(22,23),(99,99)), 0,  9) -- 14197
,( 11, E,0,0,((20,23),(21,21),( 4, 5),(22,23),(24,25),(99,99)), 0,  9) -- 14198
,( 11, E,0,0,((22,25),(23,23),( 6, 7),(24,25),(26,27),(99,99)), 0,  9) -- 14199
,( 11, E,0,0,((18,21),(18,19),( 1, 1),(20,20),(21,21),(99,99)), 0,  9) -- 14200
,( 11, E,0,0,((20,23),(20,21),( 3, 3),(22,22),(23,23),(99,99)), 0,  9) -- 14201
,( 11, E,0,0,((22,25),(22,23),( 5, 5),(24,24),(25,25),(99,99)), 0,  9) -- 14202
,( 11, E,0,0,((24,27),(24,25),( 7, 7),(26,26),(27,27),(99,99)), 0,  9) -- 14203
,( 11, E,0,0,((18,21),(16,19),( 0, 1),(16,19),(16,19),( 2, 3)), 0,  8) -- 14204
,( 11, E,0,0,((20,23),(18,21),( 2, 3),(18,21),(18,21),( 4, 5)), 0,  8) -- 14205
,( 11, E,0,0,((22,25),(20,23),( 4, 5),(20,23),(20,23),( 6, 7)), 0,  8) -- 14206
,( 11, E,0,0,((24,27),(22,25),( 6, 7),(22,25),(22,25),( 8, 9)), 0,  8) -- 14207
,( 11, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(22,25),(12,15)), 0,  8) -- 14208
,( 11, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(24,27),(14,17)), 0,  8) -- 14209
,( 11, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(26,29),(16,19)), 0,  8) -- 14210
,( 11, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(28,31),(18,21)), 0,  8) -- 14211
,( 11, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(18,21),( 6, 9)), 0,  8) -- 14212
,( 11, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(20,23),( 8,11)), 0,  8) -- 14213
,( 11, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(22,25),(10,13)), 0,  8) -- 14214
,( 11, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(24,27),(12,15)), 0,  8) -- 14215
,( 11, E,0,0,((20,23),(18,21),( 1, 1),(18,21),(20,23),( 6, 9)), 0,  8) -- 14216
,( 11, E,0,0,((22,25),(20,23),( 3, 3),(20,23),(22,25),( 8,11)), 0,  8) -- 14217
,( 11, E,0,0,((24,27),(22,25),( 5, 5),(22,25),(24,27),(10,13)), 0,  8) -- 14218
,( 11, E,0,0,((26,29),(24,27),( 7, 7),(24,27),(26,29),(12,15)), 0,  8) -- 14219
,( 11, E,0,0,((20,23),(18,21),( 0, 1),(16,19),(14,17),(99,99)), 0,  8) -- 14220
,( 11, E,0,0,((22,25),(20,23),( 2, 3),(18,21),(16,19),(99,99)), 0,  8) -- 14221
,( 11, E,0,0,((24,27),(22,25),( 4, 5),(20,23),(18,21),(99,99)), 0,  8) -- 14222
,( 11, E,0,0,((26,29),(24,27),( 6, 7),(22,25),(20,23),(99,99)), 0,  8) -- 14223
,( 11, E,0,0,((16,19),(16,19),( 0, 1),(18,21),(14,17),(99,99)), 0,  7) -- 14224
,( 11, E,0,0,((18,21),(18,21),( 2, 3),(20,23),(16,19),(99,99)), 0,  7) -- 14225
,( 11, E,0,0,((20,23),(20,23),( 4, 5),(22,25),(18,21),(99,99)), 0,  7) -- 14226
,( 11, E,0,0,((22,25),(22,25),( 6, 7),(24,27),(20,23),(99,99)), 0,  7) -- 14227
,( 11, E,0,0,((14,15),(14,17),( 0, 1),(18,21),(20,23),(99,99)), 0,  7) -- 14228
,( 11, E,0,0,((16,17),(16,19),( 2, 3),(20,23),(22,25),(99,99)), 0,  7) -- 14229
,( 11, E,0,0,((18,19),(18,21),( 4, 5),(22,25),(24,27),(99,99)), 0,  7) -- 14230
,( 11, E,0,0,((20,21),(20,23),( 6, 7),(24,27),(26,29),(99,99)), 0,  7) -- 14231
,( 11, E,0,1,((12,15),(14,17),( 0, 1),(18,21),(99,99),(99,99)), 0,  7) -- 14232
,( 11, E,0,1,((14,17),(16,19),( 2, 3),(20,23),(99,99),(99,99)), 0,  7) -- 14233
,( 11, E,0,1,((16,19),(18,21),( 4, 5),(22,25),(99,99),(99,99)), 0,  7) -- 14234
,( 11, E,0,1,((18,21),(20,23),( 6, 7),(24,27),(99,99),(99,99)), 0,  7) -- 14235
,( 11, E,0,1,((14,17),(16,19),( 0, 1),(16,17),(99,99),(99,99)), 0,  7) -- 14236
,( 11, E,0,1,((16,19),(18,21),( 2, 3),(18,19),(99,99),(99,99)), 0,  7) -- 14237
,( 11, E,0,1,((18,21),(20,23),( 4, 5),(20,21),(99,99),(99,99)), 0,  7) -- 14238
,( 11, E,0,1,((20,23),(22,25),( 6, 7),(22,23),(99,99),(99,99)), 0,  7) -- 14239
,( 11, E,0,1,((18,21),(18,21),( 0, 1),(12,15),(99,99),(99,99)), 0,  6) -- 14240
,( 11, E,0,1,((20,23),(20,23),( 2, 3),(14,17),(99,99),(99,99)), 0,  6) -- 14241
,( 11, E,0,1,((22,25),(22,25),( 4, 5),(16,19),(99,99),(99,99)), 0,  6) -- 14242
,( 11, E,0,1,((24,27),(24,27),( 6, 7),(18,21),(99,99),(99,99)), 0,  6) -- 14243
,( 11, E,0,1,(( 8,11),(12,15),( 0, 1),(18,21),(99,99),(99,99)), 0,  6) -- 14244
,( 11, E,0,1,((10,13),(14,17),( 2, 3),(20,23),(99,99),(99,99)), 0,  6) -- 14245
,( 11, E,0,1,((12,15),(16,19),( 4, 5),(22,25),(99,99),(99,99)), 0,  6) -- 14246
,( 11, E,0,1,((14,17),(18,21),( 6, 7),(24,27),(99,99),(99,99)), 0,  6) -- 14247
,( 11, E,0,1,((20,23),(20,23),( 0, 1),(10,13),(99,99),(99,99)), 0,  5) -- 14248
,( 11, E,0,1,((22,25),(22,25),( 2, 3),(12,15),(99,99),(99,99)), 0,  5) -- 14249
,( 11, E,0,1,((24,27),(24,27),( 4, 5),(14,17),(99,99),(99,99)), 0,  5) -- 14250
,( 11, E,0,1,((26,29),(26,29),( 6, 7),(16,19),(99,99),(99,99)), 0,  5) -- 14251
  );
end RPC_PAC_patt;